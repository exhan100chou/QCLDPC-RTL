module LDPCg5p16codec(
                         RESET_N,CLK,
                         start_encode,
                         data_in_tx,
                         data_in,
                         start_ldpc,start_Ldata,
                         maxiter,
                         encode_fin,
                         parity_r,
                         hb_count,
                         addr_count,
                         hardbit,
                         enga_en,dec_fin,dec_fail,hb_vlid,
                         ch_counta,ch_countb);
input        RESET_N,CLK;
input        start_encode,start_ldpc,start_Ldata;
input  [4:0] maxiter;
input  [15:0] data_in_tx;
input  [47:0] data_in;
output [3:0]  hb_count;
output [3:0] addr_count;
output [15:0] hardbit,parity_r;
output        encode_fin,enga_en,dec_fin,dec_fail,hb_vlid;
output [12:0] ch_counta,ch_countb;
wire       encode_fin;
wire [15:0] parity_r;
wire [3:0]  hb_count;
wire [3:0] addr_count;
wire [15:0] hardbit;
wire        enga_en,dec_fin,dec_fail,hb_vlid;
wire [12:0] ch_counta,ch_countb;

LDPC_enc  LDPC_enc(
                   .RESET_N(RESET_N),.CLK(CLK),
                   .start_encode(start_encode),
                   .data_in(data_in_tx),
                   .encode_fin(encode_fin),
                   .parity_r(parity_r) );
wire [47:0] chdata=data_in;

LDPCDECg5p16v8 LDPCDECg5p16v8(
             .CLK(CLK),.RESET_N(RESET_N),.start_ldpc(start_ldpc),.start_Ldata(start_Ldata),
             .maxiter(maxiter),
             .chdata(chdata),
             .hb_count(hb_count),
             .hardbit(hardbit),
             .enga_en(enga_en),.dec_fin(dec_fin),.dec_fail(dec_fail),.hb_vlid(hb_vlid),
             .ch_counta(ch_counta),.ch_countb(ch_countb),.addr_count(addr_count));

endmodule
module LDPC_enc(
                RESET_N,CLK,
                start_encode,
                data_in,
                encode_fin,
                parity_r
                                    );
input        RESET_N,CLK;
input        start_encode;
input  [15:0] data_in;
output       encode_fin;
output [15:0] parity_r;
parameter    cir_lt1  =256'b0100100110110111001110101100001010010101100000111111111011010001111101111001001100110101110110100000001011000000111110100000001111010010100011010001010101111110101111101011000001110011000001001000010100011110100111011000001001001100101000101000110010000110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt2  =256'b0001001010000010111111001000011100010000011011000010011101010010110001011111010011100010111011011010111001011010101111100110110101101110001011000111011111101010111111011101100000100010100001001101011000011010101110110000010110010001010100101000111011101000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt3  =256'b0110000001101101111111110001100001101000110111110011110110000100100011100000000101000111101011000001110001001110111111011111010011111010101110110011100101001011101111100101000010110101111011001100000111101001001001000001110100001000011001111110000000101110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt4  =256'b1011101101011000001110010101110111101101001100001110010000000111101111000110011010010000100110111011000011010100101110011001101001000110000110100101101111011111111111010011100011100100011011001001001011101101000000101001101011010101100101111110001001000000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt5  =256'b0011001001101101011101001111100110111011001000000101010110010010011111011110110000001111111101010101001111011001101011010010010001001000100111011110110100101011110101011100010111010000110001101011000111110100000111011010010010111111000000110000110000010000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt6  =256'b0010010111101101001010110001101111001000011100111001100001011100110000101100011101001111000101011111001001011010100101001000111010011111111000110111100100000000100100000001101101101110101001101101110101001111100011101100000110100100101110101100110000011010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt7  =256'b1001111110101000110100100110111100100000101110000110111101101111000101100110010000001100110011000100100001101010110111100101110100001111100110011000001100101011110010011001001011100101100010001100111010000100001000011000101110001001111001101111101111001000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt8  =256'b0000100000101000100011011000110101010011111010111010001010100001101010010100111101001100001011001110100111101001111001111111011111011000111001110001011100000000100011000100110001011011111010001010001000111111101100101110111010010010010111110011101111000010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt9  =256'b0111110011111011011001111111010100001110101110110111100111011000100000011001001100010010010111110111110110101010111101001001111000000111101100011101111000011000100010100111101000001111100100011101110111110001101101010111101010100100010111110100111000101010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt10 =256'b1011001101110111010011011110101110101000101101100101101000111000110001101101001011011101111110011011000111100110001010001111001110111110010011110110000001101101011101110010001011100001110010101010011110000000101100001101100010101010110110001011110011111000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt11 =256'b0010001100000000000010111111001110100110001001101011101101001111100100001011011110110000101000101011101100000110101111101100011010001001011100111111100000010100110000001011110110001111000111011000010010101101101000111111111111111001101110101011001001111000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt12 =256'b0110110010001100001000011110110100000000001010111001100010101111110101111111011001111111000001000111011101001010011000101010101100110000100011010100011001100001001111011110010101100001010001101111111011011100101001100101110111110111001111010100000010101010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt13 =256'b0001100101010011011001001111010001110101001101010000010011000101100010101100010111100101010101110111000011001001101101100101101110010001110010010011010101010100100111001101001100000001000111100101111110010001010110110000100001010110011010010000110001110100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt14 =256'b0001000000111000100111110011001000111110100101100111001010001111011010111010000100101011010001100110010000000011100010110100100011100110100100010100101010111011101000110010010001000110101010010110100100011100110010100110101000101011111101111010110100110100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt15 =256'b1101100101011001111100011100011010110100111110111011010011111111110001011101001101010101101010101101100011101101100110011100110001101010000100011101011111110101001101011001100111010100111010001010001110011110111110001001110010001101010010101100100001001010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt16 =256'b0101000000110010000010100000000011111111010110001100001010110101001001001011011110011011101110111100110000100111101001001101111100011101010010011010100000011010000010100110111010010011010111111001010100010011011010011111111011110000110101000110100100001010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt17 =256'b1010001110111110001001110010100101111000100101111010111100101110111000001001011100010001100110111111100100100011100010111010111000111010010001000011010000001011010001111010001010100100010000100110101110001000111010010011010110001011111100100101000101100100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt18 =256'b1011111010000100000100101000000101000010010001011101101101001011001000100011010000001110100111011010011111110010111010010011011110010000000100000111010011001101000110001101111100010011010101001011100011110100101010110111010000000011010011100110111111011110;                                                                                                                                                   
parameter    cir_lt19 =256'b1010100100000001111110010010100011110110011010010001100010110100110001110101100111110110111010100111000010010000000111111100111010011011111101111010000101111100101101000100001000101101100011010000011101100110010110110111011110110100011011110010000100011100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt20 =256'b0011010000111011110011001000000011001100101110110110110011010001000001011111101011101001111011000010111001000001011111010101011100110001101000111110000110111010111010110011111110011010100110111101010000011010000110010011011000111100110100110001111110100110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt21 =256'b0000011011000100000011100001101111010111000110111010100000011110100001010001010000011111101110010000000010010010111101010111111101011110000000111010110101110001110001101011111000101100111101001011110100000101010001001101101111011100101101000101000100000000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt22 =256'b0011110000010111001101110010101101111011110001111010010110101001110101010011010010101001110000100010011101011101100111010011111011110011011001011110000010101011111110110110101111000010001011110011110000100001101100011001111100110101011000000010111100010000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt23 =256'b1111101100001010000100100101111010111010000010101011001010111000111011000001111010111001001100011100110110010001010001000000001111010001001100010101011011111010011101100010110010111000010001000101001000000111010010001001011011001001110110001001001111101110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt24 =256'b0100000111011001001010110110111000010110110101101011111100001111101111000011111000001111010010101110101001011110001011000100001001111100010101110001101100100000010010111111100101010110100111111101001100100011101111011101001000100000000011001110110111111110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt25 =256'b0001101001100010000101000010010111110111110000010011111111101100101111110000011000000001100011101001001100110010111111101000110011101001000010100001110110111111001000010110000000100010001001111011101100010010000000110010111001111111011001100001001000111010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt26 =256'b1100100111010001000000011011111100100010011000111001001110100011000101101110110100000011111100001101110101110101111010000001010111100101010001101110111101001010011001011010010001111011101111111110001100111101110110100101001000010100110000101110100011000010;                                                                                                                                                
parameter    cir_lt27 =256'b1001100100110101000111010010010000001010111111000000010010011010110101010001111010101101100000100001011100001100011001111110011001011001010011110110010011111000000011000001111000101000010010110000100100101111010010100010110101111000000101010001011011110100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt28 =256'b1100101010000110000010001011111011011111010111101010100011010101011111001111010110101111111111000101100101001011011100010111111101010101000000111001011000001101010010001101101001110001110100110101000100000000100100110101000100010011101100011110110000001100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt29 =256'b1010011001111101110101001111000110001111111001000001101010000111111000100100000011000110110110111010111111101000110000010101101010011010010100010011111110001101101000110001001011101111100011111001100001100010100011001100100010100011101010111010010000010110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt30 =256'b1001111011000111000000110000111011011100100000101000000110000111000110000111000000001001100100010100111101110110111001100111110110010100110011111000101111010011010101000111100101011011000000001010011100101001000011111011100001110100010111100111001001000010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt31 =256'b0000111101100110010001001111000100010111000010101110001101001001101100111001000110001100001100110011011001110011101110100000100001000101101001100010011101011000100011010011000110011111011110001111010101110001011100011001010100010111010000101010000100010010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt32 =256'b1011011111011100100100110000111001000100011011000111100001001001010010011010000101000011011110011101011011101101100111010010111101001011001110001001001100000110011110100101101000101011111101111100101000111010111100101110010111000000101101110111011101000110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt33 =256'b0011010011001111101101011100110001010110111011111101001001100001000011110010111111001011000011111101111111011011000001111001111101111010100100011000010001111111000110000101101011000001110110011011000100100001100010111111101100000110110010110010000001011010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt34 =256'b0101001100010100111100011100100011101001111001100111001101010001001011001001010110101000001001101001100011101110101000111110011100110001101010101000000111100110110011000101111100101101111101100111001011011110000100101010100011001010111110010011100000001110;           
parameter    cir_lt35 =256'b0110000100111010001000001010011111001100001101000010111101011011000111000001110110010001010110100110001110001001111111101001010000101001000101110010110010010000000010011101101001001100000010110001110101110001000000100110010110011000011010100101001000010000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt36 =256'b1000011011100001011001001010001101110011001111011000111001101011001111111010011111110010011100110010010010111100010110101110110001100010001011000010100100001001110111011101111110100000001001001101111010001110100110110011011001010100010110000100101001000100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt37 =256'b0010011011110101111111011000101011010010100100001001001110011001111011011111110000000011011110110001001000100001111011111101100100111110010111111011000110010110010001011100000110001100010100010000010100111010010011010011110110011100111011011101111100101010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt38 =256'b0001101101100011000101101001111000001001100011000100010000000100001001000000111110110010000100100010100110101011001001110100100111100101000100001011100101111011100000010110001000101110110011111001010011000001000001001011111010101010111000011001010010100100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt39 =256'b1100111100011001001111101001011001001110100000110000110110111001001101110011001001010100100000011000110011100110110010100100000101100001000110000010011110001011101010101001111101110001010010111100100110110101011000010101001111111011101101111010110011010010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt40 =256'b0111001010001111110101011000001010010101100111111101101000100100111111101100000111100101111010001011011101101100000000101101000110111010010101110010111101100110011011100011110011010011110101010101100001001110001010001101000011001101101110111110011101011100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt41 =256'b0101000110100010011011010010111100100011110100011101101000010110001101110010001001000000010101000001110101010111111011100101100010001111100011010001100100110100111101001110010011100001010011100101110011100001001110101010010101000010010010010111110110111110;                                                                                                                                                   
parameter    cir_lt42 =256'b1011101100010011100100101000010011110010010011110010001000111110000101010000110001000001111001111010110001111100000010011110101001100000100100101101100111100101110011001100100110010000000110100011101011001101001001110010011011100000011000101101111111001100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt43 =256'b0010000000011010000011000111101101111101100110110000100001101010011110110111011100001101110001100000100100100010110010010011100010101111100011111010011001110000110101100100000100010110000000010011110001001110010010000010010011010011110011000111001011111100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt44 =256'b0100101010101011111100111101000010101100000001011111000001000010010110010101100100001100011101011011100000001001001011101000101001000000100100000110011010100001111011100110110001100111010101010101101001100010010101011010011101110001111001111101000010001110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt45 =256'b1100000011010111101010011110111100000001100101110011100010101010011001110111100000011010001100010100001000111101001101010001100010010100111100000101001100111011011011000010011010010001111000011001001101010110100100101011101100100001011010101100100011101100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt46 =256'b0110011010111010111000101111010111111000010001000011010110010100010011101001011101110110011010000001101000100000001001101111100000011000111100010001011111100111000001010000001101011001010011000011110000001011101111110110000010100111110011100010101100011100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt47 =256'b0011010000011111111110100010110000110011011110001011101101110110100111111101100011111011111010100010010011101011010011001100100000111100011000001100111011111011111101011111110111100000010101111001001100000011011111110100110000011100011111011010011010010110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt48 =256'b0001001001110010101100010011011011001010101010111011011001001000101101100011011110010111101100110111110011110110010111110010100010110000011000011000101000100111100111001101100000101000111110100011110001011110010100101001011110011010110110010100010101100110;         
parameter    cir_lt49 =256'b0010110000010111000000000010110111011001100100111100000001111011110001110111111011101011110011010010010111000100010100100111011100101100101001001011100011011000001111100001001110111010111101101110010001011110010011000010100001110100011111000011100111101100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt50 =256'b1010011011100011100010011011100010101000001011011011100000000100010000011110011000001011111011010111100011111111010000101001111011011111111101001000001111000001011101111101110111111001110100011001010010000100000101110011010001111100110000100110001100011000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt51 =256'b1010010010111001000001111001101001110101101001000000011001001110010100011101111100000101101010001010001101111010101111000111100001101011001010010100001110111010100110111110010110110011000100100111000001100000101011110111110001010110000001110000011000111000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt52 =256'b1010111001001101100011100000111100000100000110100111111000110001110101110100011111100101100010001111111001000001101011001001000110011000011110010111100010100011110100100010101111110000001101010000000010111010111101000110000001011110101110010101110011001100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt53 =256'b0010110111111101011111101000101000011110100110100001101000111010101010101101001101111011011110100110100110010011000000110001100101101001110110001011101010111110000001010101100100100110001100110010110001010110110100100001011111010001111011001011100101011100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt54 =256'b0111101111000010100101001010111100001010100101010100101011011000100011001111110001001110100010101001000111011000110111110001011111001011010100010000011100011000000000111010110101000010111000111110010100011000110011010011001100100010101111001011101101000100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt55 =256'b1011000000000010010101000010011010000010010011110011001001001100011110011100000000011101101110000110010110101111110101000000000010011101000000011001010011110001001011111010010000011110110010110101000100101100101101111101100011010100110000100010011111011100;                                                                                                                                                   
parameter    cir_lt56 =256'b0110011000111101101111100000001110010110010000000110001010101110010111111110111100101000010010001001110111100100000010000000111000111111100010000010100101010111001010010101000001111010000110111001100001100010101010001111110000100111100100100010010111000100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt57 =256'b0101100010011011001010011000100110110100101110011100000011110010101010111111000011000011010010000001110101100010001111100100110111100100110111110111111000110111101111001001101110101011110001100000101011110101010010010001110011111110101010100001101001100110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt58 =256'b0011111010011011000100101011100001000000000100010011101101010000010011100001010011000111011110011100000110000010100011101000111011000011111010110111101001110111101111010111101111101010101010101110101010111100101101111101010111111000000111110001000100000010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt59 =256'b1100111011010111111110011010011100000110100101101110111110001100111010111111000011101111111000101011111100000111111111001010000011101011001010101101101011011111011100100110110011100110001000000110100110100010000110101011110000000010111110000111111001101100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt60 =256'b0010100011010111110000101001011011110010001111100001010000101110000011100001010011101011110100110110001111100111010011000110001111001100000111101101111010011111011100111000110010100111010011001000100111101011111001000111010100000100010011010111010100001000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt61 =256'b1001100001011101110001111010100001001000111110111110011110000100010001111101111010111011111100011001000001111010001110100011101101100001110111011011110110011110001100000110011101001011110111000110001011010111010011101001010111100001000010100100110010110000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt62 =256'b0110001110101100111100100101100001010011100011110011001100100011010001100100011001111101101011111000001110100011110101011101111001000010110011110101001100110011011100110000001010011110100110001001111110100111110010001100010111110101101110000110001111110100;   
parameter    cir_lt63 =256'b1111011110000001100011111100110100110100001111101001111110100110010110110111011101011000000110001100000101100010001110101111101101001110011100101011000110111000111101111100011101010111101101000111010101110010011101010110100111100000000100000000001100001110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt64 =256'b1000110001110000101110100011110100101111010010100100101100000001010110101110111110011110010001101101001010111011110101010001111001101101011000000101111100010101101101001010001010000010111100001000100000000010111100110011100111110100101000100010110001001010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt65 =256'b1000101100001010100001001100000011001010101010110100000100101010011110010001000011000011100001010110110101110001100001100011110010110110111101101001110111010100010001110011000010010100101001111101101101111111001001100011101010010100100110000110000010111010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt66 =256'b1111011011110101101100111101111010000100011110011110000101110010000100111111000111001010110001101011110001011111001110001001100110111101100111111010111100000110111110100001001111001101010000000000000000110111100010111000000110001010000111010101111100000100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt67 =256'b1101111100011001001110001101010111110011000101010001010001110010011111011100000100011101000100000111011101000011010001010111110001011110111111000111010100101110001101101000010100000000011100010100011000010011110001100001001011000001010110100111000100101010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt68 =256'b0010001011100110000011111100101110111101110001111011010000101010000101110010000000010100010100111010011001101101111110111101100101010101100101010100011111111100100010111010011001011001100101101001110101011011011010111010100111011111110111110100111010010100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt69 =256'b0000101100111100100011101000001110111011011001101001010011000100011100010101101000110000000010001101011100000001011110011110010000011000010111111000011010110011011001110111101101011111011100001101001000111010010100001100010001110001111110111001110101100010;                                                                                                                                           
parameter    cir_lt70 =256'b1000001000000101111100100100110010100000010101011101010100011110011110100111101100111101010110110000000101110001100100101010100100111110111001010110000100000110001101110010001111101101111101101011111110101000000110111100011101111100001000011001001111101010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt71 =256'b1000100110000001010001110001110110010101101000101111111010111011111101000110100110001101101010011110101101001010010100111000111100001110000100111101011100011000100010001111000110010100100000010111111100001100100100100010011000011111001110001111111001100100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt72 =256'b1000000010111000001110111101001010001110100100011011111101100001111111110100100010000000111110100011110100111010101110001100001000101000101010010011000010101101110110001010100100100110000001110001001010011110110110010010010100010010111000101111000011101100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt73 =256'b1100001110001010111000000111111000111010001010111100000010100100001011101010011111010111000111110010010011001001001100000101111001000111111110100001110101100001100101101110111000111001000110011111000110111010110000100111101110011001011011110100101110011100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt74 =256'b1100110010001111111101001001000000010110101100001000000000011001000010111010010101110001001011010110001010101001110010001011010111101010000100011110110111000100011010110100011101111001000011100010001110011110100110001110111001011110110111001100101001011000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt75 =256'b0111000000010101010110000000111101001011101001100000110011110110010011000010010101101001001110011001011110110100001011010011110001111110101111100111010111111111111100010001111100011111000100101110110110001111011011010111000111100110000001011101110011000110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt76 =256'b1111111100010000010011001110000101100111001111010100110001001011011010010010011111001111000010111101000111010100110101011101011111010011010101011000010101011010000011001011011001011111000001010011111110101011001101111110010000100001101101100101110100000010;                                                                                                                                                                                                                                                                                        
parameter    cir_lt77 =256'b0110001010011000010000000010110011101100011010011010100011110100110010100101110110101011001010111110001000101001101100101011111110011011110001111100000110000111001010000010101101101000000100101111101001001000011011110011011011101100001011111111010110100100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt78 =256'b1111010101100001011001000010100111100111011000110100011010110100010101110011011001001011100111010001000111010110100010011100010000001111111011101111101011000100000001101100010010110000000001111011101001101010110011000100101111001110111111101011100000111100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt79 =256'b1110110001100110001010100111110001100101100100000111101110000001000001010011010010010101111111111010010100000001011010001011110000001000100110111110000000011001111101001101001000000000010000100101010110101111100101000000011010111110000110011101101100110100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt80 =256'b1111101110011111000011100111100101101110100110101001010111000001100110000101111101110101010010010101011011111110010100111100011110011100101100101101101101011010110110100011110111011000010101110001010110001101001101110111101110011100110010001001011010101100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt81 =256'b1101100001010000011000110000000100000111101101010001010010110001010000000100110010100010011101111101101011011001101100101011001110010011101110110111000111111001111001011111011110101010000100010010100111111111001100100101011100000000011100011100010101001010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt82 =256'b1101101111100111001100100100001010100010001011110000010001110100101111110011100001011001000010110101111101000010100011001010000010100111001101110010111010001001111110001001111100010110111001100111101011011101111000110110110000001010110100101111010010011100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt83 =256'b0111011011111101010100000011010001100111100011011011010001001010110110000011001011000010000010011110110101010011000100110000101000010100010001110011110101000101000011000001100101111110101001001001100111011110011000101111101011001000100001100001111010100010;                                                                                                                                                 
parameter    cir_lt84 =256'b1111010101001010000000010111011111000010000101111010010010001111001001110100011000111001011101010110100011001000001011010001100100100000110010110110001000110101000100010111000111000010010100111100101011111100101100111100000111000010001001010010111101110100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt85 =256'b0011000001100001100001000110110011100000001101110001001100100110110110001011001111001000001001110010001100111001001110111011011011011110100110001101110001100010110010101101100011010010011001010001000110001010110001100100101111001001110000010010010010011110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt86 =256'b1111110100000111001101101000000011001110011111100101001001110110000010101010111000110110011101010101111001110111110110101011011000011000101110011000010110110001100000111110110111000111100110010110100101011001010001100010101110100111011111000000101110110100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt87 =256'b0101010100001000001000011110010010110000110010101000101101000000101110111000010001111010111100111111101111010100001000010001000101000000010101100100000001010101000110101110000100111010001010000011100011010000010000000100011001110101110010111100100010111010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt88 =256'b0001100001101110100100110000100010011110100000111100101000010000011010011001100110000100101000011000011010011010110000000001000110000110011101110001100110000110010100111101010000101111110101000100000000000011110000000010011000011011011101101110011110010000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt89 =256'b0000001010101111001001001001100011100010011000110001011000000101101111111011110011111111100111101000110000100001100110110111001001100011100001100111100001010101101111000101000001101101100000000111101010111111101100011101010111100001100010100010101001111000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt90 =256'b1000010001000100011101001111000001110010000110011000101100100111110101110001101010001100001011110000000100100011110010001001110111101000011100101001011110000011101111101001101101101110010110010011111111001100011010101111000010011001001100111001110100010010;                                                                                                                                                                                                                                                                                               
parameter    cir_lt91 =256'b1100101001111000100100001001000010101001100011100111100011001111000100111111110000100001100110001101000111101010000011001101000111011100110001101110001100111110101000110110101100110011110010011110101000001100101100011001110101010010011000111110000010101010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt92 =256'b1100110010010011110000001111100000111001111101001110010111101101011110110101101001010010001010010101110011101000010111110011111001010111001100100000110011101000101000011010000000110000000100001010111101111111011010101011100000101010110110100101011111000000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt93 =256'b0110111000110010000010000110011011111101011011010101010011011010110100011001001010111111110111101000100111000100011110100001001100001101010100011111110100011011001111001011000111011000110000010110010001110100010001011000010110111011011110000000101000101000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt94 =256'b0100110010100101011101101011011100110010101100010000111101110110110011101011011111111000011010101100010111011011111011111000010100111000011001111100110001101110111111100110100101010101000000110101111011110010001100100100000011011001101100010101000101000110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt95 =256'b0001100111100010111100100011101000111100111100010000000010000011010111001001010111111011111000000101100110110010011111100011010001000111010001110000011000011001000101100010000100110110111001101011001110110101010001100011111101101101111111101001101010000000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt96 =256'b1011101101110101100011001110101111110011001011010101101100101111010000111011000010111100010101000001010110101101111010111010001001110010011100010011011101101100110101001111100110111011001001001000100100110011001100011111101000001111001101111100000111101110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt97 =256'b1100111101010000101011010110100010100000100110101010100011111001011100100101000101111011110110001011010110011001101110000010110110111000100101011111010101110010001100011000101011101001001110110010000100011000010101100000100100100100110010000000101000000010;                                                                                                                                               
parameter    cir_lt98 =256'b1000010001011110111011110110111001101110010011111000001000010100101011101101010111001110100000101000110100010111100000001110111001111101111000110011000010100100100100110110001001100101101111111011100111011100010000011010001001100011000100000101000101000100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt99 =256'b0101101000101000010111000010000100001101010011011100111000110000110010101000010001001011010011010100010001101010100110001011101011111101000100100011111100011111000111100111000100110001000010110000010011111111010101000101100001010111001011010100101111100000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt100=256'b1001000100100110000111100010011111000011100110001110010011011101000101100000000011111110000101110111110011100100101000000111100100111000011001001111101011001001101111001001100110111101100011111001110000111011010000111111001100010000111101010001000010100110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt101=256'b1001101111100110001100110011101000000011111000010000101010000101111100110110100000011110100000110000001111110010010010101010111110011101101010011110101011011000110011110011100101101010001100011001010000101111111101101000001010010000100011011001101100100010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt102=256'b1101011100111010000101000010111011101101011100001001111110111110001001100010001001110110000111101010010110111111011110111000101110011111010000010011010111110010111010110001001100000110110101001000010101000011110111010000110011010100101001110011000100010010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt103=256'b0011000001010000011111000100101100010101010101110100111111001000011011110111100010010110100110101011011001011101110011100001010000011011001010111100100011010011101010001101111100010001101011101011111100100101001100111001101100001100110111000011001000111110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt104=256'b1111110010001100010110110101111111111011110001101101101011110011101110100011001011111110000001110001000000010000111111110011000000011001110000110001011111111001100011001111010101111101010010111010111001001001000110000001010101001000111101101001100000001110;  
parameter    cir_lt105=256'b1110011110111011010001111101010001001011101011011001000111101101111011100000101010011001010000110101010010010010010110111001110011001111111111110000001101111011111110000111001111110001000010101000011100100101010111000111011000111011001100011011111011111100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt106=256'b0010000111010010011111010110001100101010110011000111010110100100110100100100001100100001001000010000001110001010100011010001100010000111110010101101000111000110010010100110000101011111100110001001000100101001110000100111011000010011000100011101111001001100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt107=256'b1110001110000111011101001110111000010000100110001111100101011100011000001000001111010001110010110101110001111111100000010101110001001100100100110111111011011001110100011011001001111010010010101001010001100110001101111100110000000110101000000111110101100110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt108=256'b1010010111101110010011100101100101110001111110010001110100010101010111001100101001101001101010010000101101100111010101111101100000000100101001101010110001100100011000111010000011010100110110001000001001101010101010011100110000101110100000000001110111010110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt109=256'b0011101011011101110001111110011111111010001010100110001011010001001101100100100011001111111001001111101001101001101011010100110001010011010111011110001001011110000110111000000001111010100001000111011111100111001001010101011110110010110000110100101001111100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt110=256'b1101000110001010100100111101110111111001000111110010100010000111011010100001111100100011110011010001101100101010001100011011011100011010000110101010011100101010001011110001101010101111100111111110111111000111010000100001110011000010000010010110001011011010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt111=256'b1000111001111010011100000111100101100010010110111011110011010111100100011001000101100110101000001101111100011100111110001001101011111101110001111111101111100010001110001001010111101001110100010001110011101100010100111101011011101000101010101111000011010110;  
parameter    cir_lt112=256'b1110010100101101001001000100001101100001011011101111011010000001110011011100011010001010100010010011111001011111011001000110000110110100100000001011111010010110000011000000111100111100110010101000010011001100001101001001110110011000011000001101100001110000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt113=256'b1011010101000011011110011111001110000011111100000111011001000101110111011001100110000101001011101011010110010100101011100010000100100010011111011100111011111100010010010000010000001011010101101010010100110011100010111000010110000010011000001100001011000110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt114=256'b1111000001110001001001010101010000100111000111100110000010111000011110001000011100111101011111010101001000111011111101001111111011110000010010001111100101110100100101011011000100001110000110111100011001001111010100011110001011011011000110000110111001011110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt115=256'b0000101001001100001001111011101001011000010110001011000101111111101011000000001011011000010010011000010011101011110101000001110101010100100001010011010100011000100100110011001100001100001101011100101101010110100000111011100000001010101100010010111011011000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt116=256'b1100111101111110011110110001110111111100101101101010011110000010000010010001110001100000000110100110001101000100100011101100001010000110101100000000001010010000010011111000011000001001011110001010100000101010010110011101111101010011110010011000001001000000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt117=256'b0110100111110100000010100001100111111000001100101110010110110110111111111000101110010000000110000001101010000011110101101001001110001110011110011100100100101010101010100111111011110011010101001101010111000011100011110011111001000100001111000100110010011010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt118=256'b0000000011111011100010010010101100001000101000000100100111000111001011111101100001011101010010001011000000110110000101101001010101111000000010010000011111001101010010000101001111100111100011110010101111101010111100010110100111001010101000010111001001101010; 
parameter    cir_lt119=256'b0010111011011010101110100001111101100111011111011110010110010001111110000001000000101011111011001111100000001000011011000010001111100001000101111010000111000001011010011100111010000011011111010100000000011001001100100011010100010001110001101011011101001100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt120=256'b1100011111010101001110010010110110010111111011110100100111100000001010000100001111100110101111000101001010111101101011000010010100010111011001110110111100100110100010111110001110010111101001101011111000110000010011000110001010011111010110111000100110111100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt121=256'b1011101110001110111000100101100111011110000010001100011010010101001100011101011100010100110001110000001100011111110110000010100110000001100001101000110111000101010111000100111010001110111110011101000110011000110011010001001000100111011111001111000110010000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt122=256'b1001110011001111010110001000110011101110010110101110101010001001100100101000110011101011011101010000010111110001111111000110101011111010011000111100011011110010000100011110001001100001110010001010100001110000001011011001011000001000111001100011000010000000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt123=256'b1111000100010010001101110001110011100101101000011111100000101100010111010110000001100110011111010111100110110010100001010010000011101000011101100110010110101001010100110111000100100001100101100000111110110000110110110101001111001101100100010011010101110110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt124=256'b0101011001010011100011011100100111010101111100111101010000110000111111100011101110011001110011110111111101011100101000010110001110010011100100110010111010011110000111101101110111001110101001110111011001011000001110111101011111100010000010111111010001100110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt125=256'b1111101011011000100011011010101000010100011010101100000000011111101111111000110110101011111100111110000101001010101111001100100110000000111101000101100111110011111000100110011000010010000111011101001110110110000000010101100111111111010011111101010010110100; 
parameter    cir_lt126=256'b0011110011111101011001001110100000011001010101100111110001011000100100110000001111010101111100010100011111010010101000011101010111111011111010101001011000101101100100111110110000110101001001110110001101011101010111000010100110010001010011111010101111110010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt127=256'b0110010000001100010100111101000100110000001110111001100011110010101001101100011111111000001000100110100011110000101011110011010110001010000101011010001110110001001100010010101110001001111100110110101101110010100000101001000101101100111011001000100000100000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt128=256'b0010001000101001101110101001001100111101000001110010010010110101100010100100100110000110001000001100111001101000101100100010100111110001000010110110110001101111010000001010000110101110110010011101101110011001110111111110000100000010111011001111011101100110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt129=256'b1000100011100110011011010001010001001101111111000011011100101110111100101001111111111010100101010011111011000000010100001100101101001001011101110110110000111110100000101100110010011010101111011010001000100010000101011000110101001000110000001110000100111100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt130=256'b1011110111001010100101000000111111000100010110100000101000100010001011011101100101100000110011111001101101011111101001001101100000101100101100011111000000001001001001110011001010001110100111100101000110011101010101011011110111100101000111110000100111000010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt131=256'b1100101101000001001011111110101011011110010011010111001000010000111001000001101100110110101001101001001111010111101011001011110010100001100001110100110010110110101111010111101010000110000110001011011100000001110111110000111001100000100001000100001000111110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt132=256'b0111111001101101110101101111000101010111111010110100111100011100001110110101110110101100111111000011011001001000010110001010111111000100010000011101000010000001000110001000010010010010001110110100010010111110100111110011111011001101010110111010101011000000; 
parameter    cir_lt133=256'b0100000111000010100111100001010100000110111100010111010110110100001001110100001111101001011010111100010100100010110101011000100001001101111111000100010100101001111100001111110100100100101010011011000001001101100110000110010011110001010100111001111111000010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt134=256'b0010001000010011010011101011010001100100100111001001000011000100001100100010000011001111001001110110011101010000111011101100011100101011101011011111110100000000010001110100010001011101010011001010100101100101001000000111010010111100110100000111011000101000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt135=256'b1100000001011001001010111110110011110101001011111110010101001010001001101001010001101011101010101000000111011111011001101011111101001110101101100110011000110011110011001011011010010011100101001101010011110010101010111010110000110010100111111011001100110010;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt136=256'b0010001110001000111110110100110110010111010000100000000000111010001100111111011101001101111001100010001110101101010111011111000000101000111001111101111000011010011110110000111111101010011100011100110111011010000100111011110001111111000111000101101011011000;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt137=256'b1110001100110010010010100011001011110000010101110011011000000011111110100010101110100000000011010110010010101010011001100001010110011101011110001011001000100111010000110100100000010100100111100011011110010011110111011111010011110110011000000011001100010100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt138=256'b0111110111101001001111100000000101100011110010100011010101100100010100000011110100000000011001001110101111011111000101000001110110110101001101101110100101000011100111100011011111011101100111101011011101111000000010011010111110000111111111100101000010000110;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt139=256'b0000011010011010101110111100000111010010110001000001011111100001111001110111111000001101110100110000110111000100110011111010000011110101001100111100101001010011110101001100000111100000100110010110011111011100000011001111100010100000101111001011001001111110;  
parameter    cir_lt140=256'b0001100001000001110011111111001001000001010110010001010010000110010011010110100010101101101110101000001010110001101111011010100011011101011111011001000100110111000010011011111000101001100110011110011100110111110110001010001111010001001000101101000111101100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt141=256'b0010110010110111001000110011001100100111001111000011011001000111001001000000000001101001001100101010100011000000111010101110001010010001001111000110100110011011100111101110101001100100100111100110110010001100101000111011100110001000101101100110101011111100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt142=256'b0111000011001001010000100111100101100110011011101001010011011011101101001001000001100001110000101100001001011011101101100100110000100100111000111000001000010111100011111011111101111111011111001110010011110110001010010100000010011001000011000000011111010100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt143=256'b1010110111111101001100101110111000100100000100000010011000010010100000111100101101101101000000010001000111110110101110110010000001110010001010001000101101010111001101100110010100011000110110101110101010110110000100101011000111010011001111111000011100101100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
parameter    cir_lt144=256'b0111000110000011010100111010010001100101010000101000010010001110000100110101101101100101111100010111101101101101111001111000111011000111111101110110000011011011001001110011000000000011001110000110001011001100100110000100100011000010100001011110101000000100;                                                                                                                                                                                                                                                                                                                                                                                                                                    
reg [9:0]   counter;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             
reg [1:0]   state;
reg [255:0] parity1,parity2,parity3,parity4;
reg [255:0] cir_lt_r1,cir_lt_r2,cir_lt_r3,cir_lt_r4;
reg         encode_fin;
reg [15:0]   parity_r;

wire [255:0] cir_lt_r10=(data_in[15])?cir_lt_r1:256'd0,
             cir_lt_r20=(data_in[15])?cir_lt_r2:256'd0,
             cir_lt_r30=(data_in[15])?cir_lt_r3:256'd0,
             cir_lt_r40=(data_in[15])?cir_lt_r4:256'd0,
             cir_lt_r11=(data_in[14])?{cir_lt_r1[0]  ,cir_lt_r1[255:1]}:256'd0,
             cir_lt_r21=(data_in[14])?{cir_lt_r2[0]  ,cir_lt_r2[255:1]}:256'd0,
             cir_lt_r31=(data_in[14])?{cir_lt_r3[0]  ,cir_lt_r3[255:1]}:256'd0,
             cir_lt_r41=(data_in[14])?{cir_lt_r4[0]  ,cir_lt_r4[255:1]}:256'd0,
             cir_lt_r12=(data_in[13])?{cir_lt_r1[1:0],cir_lt_r1[255:2]}:256'd0,
             cir_lt_r22=(data_in[13])?{cir_lt_r2[1:0],cir_lt_r2[255:2]}:256'd0,
             cir_lt_r32=(data_in[13])?{cir_lt_r3[1:0],cir_lt_r3[255:2]}:256'd0,
             cir_lt_r42=(data_in[13])?{cir_lt_r4[1:0],cir_lt_r4[255:2]}:256'd0,
             cir_lt_r13=(data_in[12])?{cir_lt_r1[2:0],cir_lt_r1[255:3]}:256'd0,
             cir_lt_r23=(data_in[12])?{cir_lt_r2[2:0],cir_lt_r2[255:3]}:256'd0,
             cir_lt_r33=(data_in[12])?{cir_lt_r3[2:0],cir_lt_r3[255:3]}:256'd0,
             cir_lt_r43=(data_in[12])?{cir_lt_r4[2:0],cir_lt_r4[255:3]}:256'd0,
             cir_lt_r14=(data_in[11])?{cir_lt_r1[3:0],cir_lt_r1[255:4]}:256'd0,
             cir_lt_r24=(data_in[11])?{cir_lt_r2[3:0],cir_lt_r2[255:4]}:256'd0,
             cir_lt_r34=(data_in[11])?{cir_lt_r3[3:0],cir_lt_r3[255:4]}:256'd0,
             cir_lt_r44=(data_in[11])?{cir_lt_r4[3:0],cir_lt_r4[255:4]}:256'd0,
             cir_lt_r15=(data_in[10])?{cir_lt_r1[4:0],cir_lt_r1[255:5]}:256'd0,
             cir_lt_r25=(data_in[10])?{cir_lt_r2[4:0],cir_lt_r2[255:5]}:256'd0,
             cir_lt_r35=(data_in[10])?{cir_lt_r3[4:0],cir_lt_r3[255:5]}:256'd0,
             cir_lt_r45=(data_in[10])?{cir_lt_r4[4:0],cir_lt_r4[255:5]}:256'd0,
             cir_lt_r16=(data_in[9])?{cir_lt_r1[5:0],cir_lt_r1[255:6]}:256'd0,
             cir_lt_r26=(data_in[9])?{cir_lt_r2[5:0],cir_lt_r2[255:6]}:256'd0,
             cir_lt_r36=(data_in[9])?{cir_lt_r3[5:0],cir_lt_r3[255:6]}:256'd0,
             cir_lt_r46=(data_in[9])?{cir_lt_r4[5:0],cir_lt_r4[255:6]}:256'd0,
             cir_lt_r17=(data_in[8])?{cir_lt_r1[6:0],cir_lt_r1[255:7]}:256'd0,
             cir_lt_r27=(data_in[8])?{cir_lt_r2[6:0],cir_lt_r2[255:7]}:256'd0,
             cir_lt_r37=(data_in[8])?{cir_lt_r3[6:0],cir_lt_r3[255:7]}:256'd0,
             cir_lt_r47=(data_in[8])?{cir_lt_r4[6:0],cir_lt_r4[255:7]}:256'd0,
             cir_lt_r18 =(data_in[7])?{cir_lt_r1[7:0],cir_lt_r1[255:8]}:256'd0,
             cir_lt_r28 =(data_in[7])?{cir_lt_r2[7:0],cir_lt_r2[255:8]}:256'd0,
             cir_lt_r38 =(data_in[7])?{cir_lt_r3[7:0],cir_lt_r3[255:8]}:256'd0,
             cir_lt_r48 =(data_in[7])?{cir_lt_r4[7:0],cir_lt_r4[255:8]}:256'd0,
             cir_lt_r19 =(data_in[6])?{cir_lt_r1[8:0],cir_lt_r1[255:9]}:256'd0,
             cir_lt_r29 =(data_in[6])?{cir_lt_r2[8:0],cir_lt_r2[255:9]}:256'd0,
             cir_lt_r39 =(data_in[6])?{cir_lt_r3[8:0],cir_lt_r3[255:9]}:256'd0,
             cir_lt_r49 =(data_in[6])?{cir_lt_r4[8:0],cir_lt_r4[255:9]}:256'd0,
             cir_lt_r110=(data_in[5])?{cir_lt_r1[9:0],cir_lt_r1[255:10]}:256'd0,
             cir_lt_r210=(data_in[5])?{cir_lt_r2[9:0],cir_lt_r2[255:10]}:256'd0,
             cir_lt_r310=(data_in[5])?{cir_lt_r3[9:0],cir_lt_r3[255:10]}:256'd0,
             cir_lt_r410=(data_in[5])?{cir_lt_r4[9:0],cir_lt_r4[255:10]}:256'd0,
             cir_lt_r111=(data_in[4])?{cir_lt_r1[10:0],cir_lt_r1[255:11]}:256'd0,
             cir_lt_r211=(data_in[4])?{cir_lt_r2[10:0],cir_lt_r2[255:11]}:256'd0,
             cir_lt_r311=(data_in[4])?{cir_lt_r3[10:0],cir_lt_r3[255:11]}:256'd0,
             cir_lt_r411=(data_in[4])?{cir_lt_r4[10:0],cir_lt_r4[255:11]}:256'd0,
             cir_lt_r112=(data_in[3])?{cir_lt_r1[11:0],cir_lt_r1[255:12]}:256'd0,
             cir_lt_r212=(data_in[3])?{cir_lt_r2[11:0],cir_lt_r2[255:12]}:256'd0,
             cir_lt_r312=(data_in[3])?{cir_lt_r3[11:0],cir_lt_r3[255:12]}:256'd0,
             cir_lt_r412=(data_in[3])?{cir_lt_r4[11:0],cir_lt_r4[255:12]}:256'd0,
             cir_lt_r113=(data_in[2])?{cir_lt_r1[12:0],cir_lt_r1[255:13]}:256'd0,
             cir_lt_r213=(data_in[2])?{cir_lt_r2[12:0],cir_lt_r2[255:13]}:256'd0,
             cir_lt_r313=(data_in[2])?{cir_lt_r3[12:0],cir_lt_r3[255:13]}:256'd0,
             cir_lt_r413=(data_in[2])?{cir_lt_r4[12:0],cir_lt_r4[255:13]}:256'd0,
             cir_lt_r114=(data_in[1])?{cir_lt_r1[13:0],cir_lt_r1[255:14]}:256'd0,
             cir_lt_r214=(data_in[1])?{cir_lt_r2[13:0],cir_lt_r2[255:14]}:256'd0,
             cir_lt_r314=(data_in[1])?{cir_lt_r3[13:0],cir_lt_r3[255:14]}:256'd0,
             cir_lt_r414=(data_in[1])?{cir_lt_r4[13:0],cir_lt_r4[255:14]}:256'd0,
             cir_lt_r115=(data_in[0])?{cir_lt_r1[14:0],cir_lt_r1[255:15]}:256'd0,
             cir_lt_r215=(data_in[0])?{cir_lt_r2[14:0],cir_lt_r2[255:15]}:256'd0,
             cir_lt_r315=(data_in[0])?{cir_lt_r3[14:0],cir_lt_r3[255:15]}:256'd0,
             cir_lt_r415=(data_in[0])?{cir_lt_r4[14:0],cir_lt_r4[255:15]}:256'd0;
parameter idle=2'b00,encode=2'b01,dataout=2'b10;
always @(*)
begin
  case(counter)
    10'd0  :parity_r=parity1[255:240];
    10'd1  :parity_r=parity1[239:224];
    10'd2  :parity_r=parity1[223:208];
    10'd3  :parity_r=parity1[207:192];
    10'd4  :parity_r=parity1[191:176];
    10'd5  :parity_r=parity1[175:160];
   10'd6  :parity_r=parity1[159:144];
    10'd7  :parity_r=parity1[143:128];
    10'd8  :parity_r=parity1[127:112];
    10'd9  :parity_r=parity1[111: 96];
    10'd10 :parity_r=parity1[ 95: 80];
    10'd11 :parity_r=parity1[ 79: 64];
    10'd12 :parity_r=parity1[ 63: 48];
    10'd13 :parity_r=parity1[ 47: 32];
    10'd14 :parity_r=parity1[ 31: 16];
    10'd15 :parity_r=parity1[ 15:  0];
    10'd16 :parity_r=parity2[255:240];
    10'd17 :parity_r=parity2[239:224];
    10'd18 :parity_r=parity2[223:208];
    10'd19 :parity_r=parity2[207:192];
    10'd20 :parity_r=parity2[191:176];
    10'd21 :parity_r=parity2[175:160];
    10'd22 :parity_r=parity2[159:144];
    10'd23 :parity_r=parity2[143:128];
    10'd24 :parity_r=parity2[127:112];
    10'd25 :parity_r=parity2[111: 96];
    10'd26 :parity_r=parity2[ 95: 80];
    10'd27 :parity_r=parity2[ 79: 64];
    10'd28 :parity_r=parity2[ 63: 48];
    10'd29 :parity_r=parity2[ 47: 32];
    10'd30 :parity_r=parity2[ 31: 16];
    10'd31 :parity_r=parity2[ 15:  0];
    10'd32 :parity_r=parity3[255:240];
    10'd33 :parity_r=parity3[239:224];
    10'd34 :parity_r=parity3[223:208];
    10'd35 :parity_r=parity3[207:192];
    10'd36 :parity_r=parity3[191:176];
    10'd37 :parity_r=parity3[175:160];
    10'd38 :parity_r=parity3[159:144];
    10'd39 :parity_r=parity3[143:128];
    10'd40 :parity_r=parity3[127:112];
    10'd41 :parity_r=parity3[111: 96];
    10'd42 :parity_r=parity3[ 95: 80];
    10'd43 :parity_r=parity3[ 79: 64];
    10'd44 :parity_r=parity3[ 63: 48];
    10'd45 :parity_r=parity3[ 47: 32];
    10'd46 :parity_r=parity3[ 31: 16];
    10'd47 :parity_r=parity3[ 15:  0];
    10'd48 :parity_r=parity4[255:240];
    10'd49 :parity_r=parity4[239:224];
    10'd50 :parity_r=parity4[223:208];
    10'd51 :parity_r=parity4[207:192];
    10'd52 :parity_r=parity4[191:176];
    10'd53 :parity_r=parity4[175:160];
    10'd54 :parity_r=parity4[159:144];
    10'd55 :parity_r=parity4[143:128];
    10'd56 :parity_r=parity4[127:112];
    10'd57 :parity_r=parity4[111: 96];
    10'd58 :parity_r=parity4[ 95: 80];
    10'd59 :parity_r=parity4[ 79: 64];
    10'd60 :parity_r=parity4[ 63: 48];
    10'd61 :parity_r=parity4[ 47: 32];
    10'd62 :parity_r=parity4[ 31: 16];
    10'd63 :parity_r=parity4[ 15:  0];
    default:parity_r=0;
  endcase
end
always @(negedge RESET_N or posedge CLK)
begin
  if (~RESET_N)
  begin
    parity1   <=256'd0;
    parity2   <=256'd0;
    parity3   <=256'd0;
    parity4   <=256'd0;
    cir_lt_r1 <=256'd0;
    cir_lt_r2 <=256'd0;
    cir_lt_r3 <=256'd0;
    cir_lt_r4 <=256'd0;
    state     <=idle;
    counter   <=10'b0;
    encode_fin<=1;
  end
  else
  begin
    case(state)
    idle:
    begin
      parity1  <=256'd0;
      parity2  <=256'd0;
      parity3  <=256'd0;
      parity4  <=256'd0;
      cir_lt_r1<=cir_lt1;
      cir_lt_r2<=cir_lt2;
      cir_lt_r3<=cir_lt3;
      cir_lt_r4<=cir_lt4;
      state     <=(start_encode) ? encode : idle;
      counter   <=0;
      encode_fin<= ~(start_encode);
    end
    encode:
    begin
      parity1  <=parity1^cir_lt_r10^cir_lt_r11^cir_lt_r12^cir_lt_r13^cir_lt_r14^cir_lt_r15^cir_lt_r16^cir_lt_r17^cir_lt_r18^cir_lt_r19^cir_lt_r110^cir_lt_r111^cir_lt_r112^cir_lt_r113^cir_lt_r114^cir_lt_r115;
      parity2  <=parity2^cir_lt_r20^cir_lt_r21^cir_lt_r22^cir_lt_r23^cir_lt_r24^cir_lt_r25^cir_lt_r26^cir_lt_r27^cir_lt_r28^cir_lt_r29^cir_lt_r210^cir_lt_r211^cir_lt_r212^cir_lt_r213^cir_lt_r214^cir_lt_r215;
      parity3  <=parity3^cir_lt_r30^cir_lt_r31^cir_lt_r32^cir_lt_r33^cir_lt_r34^cir_lt_r35^cir_lt_r36^cir_lt_r37^cir_lt_r38^cir_lt_r39^cir_lt_r310^cir_lt_r311^cir_lt_r312^cir_lt_r313^cir_lt_r314^cir_lt_r315;
      parity4  <=parity4^cir_lt_r40^cir_lt_r41^cir_lt_r42^cir_lt_r43^cir_lt_r44^cir_lt_r45^cir_lt_r46^cir_lt_r47^cir_lt_r48^cir_lt_r49^cir_lt_r410^cir_lt_r411^cir_lt_r412^cir_lt_r413^cir_lt_r414^cir_lt_r415;
      cir_lt_r1<={cir_lt_r1[15:0],cir_lt_r1[255:16]};
      cir_lt_r2<={cir_lt_r2[15:0],cir_lt_r2[255:16]};
      cir_lt_r3<={cir_lt_r3[15:0],cir_lt_r3[255:16]};
      cir_lt_r4<={cir_lt_r4[15:0],cir_lt_r4[255:16]};
      state        <=(counter==10'd575) ? dataout : encode;
      counter      <=(counter==10'd575) ? 0       : counter+1;
      encode_fin   <=(counter==10'd575) ;
      if(counter<=10'd1023)
      begin
          if(counter==10'd575)
      begin
          if(counter==10'd575)
          begin
          cir_lt_r1<=cir_lt1;
          cir_lt_r2<=cir_lt2;
          cir_lt_r3<=cir_lt3;
          cir_lt_r4<=cir_lt4;
          end
          if(counter==10'd15)
          begin
          cir_lt_r1<=cir_lt5;
          cir_lt_r2<=cir_lt6;
          cir_lt_r3<=cir_lt7;
          cir_lt_r4<=cir_lt8;
          end
          if(counter==10'd31)
          begin
          cir_lt_r1<=cir_lt9 ;
          cir_lt_r2<=cir_lt10;
          cir_lt_r3<=cir_lt11;
          cir_lt_r4<=cir_lt12;
          end
          if(counter==10'd47)
          begin
          cir_lt_r1<=cir_lt13;
          cir_lt_r2<=cir_lt14;
          cir_lt_r3<=cir_lt15;
          cir_lt_r4<=cir_lt16;
          end
          if(counter==10'd63)
          begin
          cir_lt_r1<=cir_lt17;
          cir_lt_r2<=cir_lt18;
          cir_lt_r3<=cir_lt19;
          cir_lt_r4<=cir_lt20;
          end
          if(counter==10'd79)
          begin
          cir_lt_r1<=cir_lt21;
          cir_lt_r2<=cir_lt22;
          cir_lt_r3<=cir_lt23;
          cir_lt_r4<=cir_lt24;
          end
          if(counter==10'd95)
          begin
          cir_lt_r1<=cir_lt25;
          cir_lt_r2<=cir_lt26;
          cir_lt_r3<=cir_lt27;
          cir_lt_r4<=cir_lt28;
          end
          if(counter==10'd111)
          begin
          cir_lt_r1<=cir_lt29;
          cir_lt_r2<=cir_lt30;
          cir_lt_r3<=cir_lt31;
          cir_lt_r4<=cir_lt32;
          end
          if(counter==10'd127 )
          begin
          cir_lt_r1<=cir_lt33;
          cir_lt_r2<=cir_lt34;
          cir_lt_r3<=cir_lt35;
          cir_lt_r4<=cir_lt36;
          end
          if(counter==10'd143 )
          begin
          cir_lt_r1<=cir_lt37;
          cir_lt_r2<=cir_lt38;
          cir_lt_r3<=cir_lt39;
          cir_lt_r4<=cir_lt40;
          end
          if(counter==10'd159 )
          begin
          cir_lt_r1<=cir_lt41;
          cir_lt_r2<=cir_lt42;
          cir_lt_r3<=cir_lt43;
          cir_lt_r4<=cir_lt44;
          end
          if(counter==10'd175 )
          begin
          cir_lt_r1<=cir_lt45;
          cir_lt_r2<=cir_lt46;
          cir_lt_r3<=cir_lt47;
          cir_lt_r4<=cir_lt48;
          end
          if(counter==10'd191 )
          begin
          cir_lt_r1<=cir_lt49;
          cir_lt_r2<=cir_lt50;
          cir_lt_r3<=cir_lt51;
          cir_lt_r4<=cir_lt52;
          end
          if(counter==10'd207 )
          begin
          cir_lt_r1<=cir_lt53;
          cir_lt_r2<=cir_lt54;
          cir_lt_r3<=cir_lt55;
          cir_lt_r4<=cir_lt56;
          end
          if(counter==10'd223 )
          begin
          cir_lt_r1<=cir_lt57;
          cir_lt_r2<=cir_lt58;
          cir_lt_r3<=cir_lt59;
          cir_lt_r4<=cir_lt60;
          end
          if(counter==10'd239  )
          begin
          cir_lt_r1<=cir_lt61;
          cir_lt_r2<=cir_lt62;
          cir_lt_r3<=cir_lt63;
          cir_lt_r4<=cir_lt64;
          end
          if(counter==10'd255 )
          begin
          cir_lt_r1<=cir_lt65;
          cir_lt_r2<=cir_lt66;
          cir_lt_r3<=cir_lt67;
          cir_lt_r4<=cir_lt68;
          end
          if(counter==10'd271 )
          begin
          cir_lt_r1<=cir_lt69;
          cir_lt_r2<=cir_lt70;
          cir_lt_r3<=cir_lt71;
          cir_lt_r4<=cir_lt72;
          end
          if(counter==10'd287 )
          begin
          cir_lt_r1<=cir_lt73;
          cir_lt_r2<=cir_lt74;
          cir_lt_r3<=cir_lt75;
          cir_lt_r4<=cir_lt76;
          end
          if(counter==10'd303 )
          begin
          cir_lt_r1<=cir_lt77;
          cir_lt_r2<=cir_lt78;
          cir_lt_r3<=cir_lt79;
          cir_lt_r4<=cir_lt80;
          end
          if(counter==10'd319 )
          begin
          cir_lt_r1<=cir_lt81;
          cir_lt_r2<=cir_lt82;
          cir_lt_r3<=cir_lt83;
          cir_lt_r4<=cir_lt84;
          end
          if(counter==10'd335 )
          begin
          cir_lt_r1<=cir_lt85;
          cir_lt_r2<=cir_lt86;
          cir_lt_r3<=cir_lt87;
          cir_lt_r4<=cir_lt88;
          end
          if(counter==10'd351 )
          begin
          cir_lt_r1<=cir_lt89;
          cir_lt_r2<=cir_lt90;
          cir_lt_r3<=cir_lt91;
          cir_lt_r4<=cir_lt92;
          end
          if(counter==10'd367 )
          begin
          cir_lt_r1<=cir_lt93;
          cir_lt_r2<=cir_lt94;
          cir_lt_r3<=cir_lt95;
          cir_lt_r4<=cir_lt96;
          end
          if(counter==10'd383 )
          begin
          cir_lt_r1<=cir_lt97 ;
          cir_lt_r2<=cir_lt98 ;
          cir_lt_r3<=cir_lt99 ;
          cir_lt_r4<=cir_lt100;
          end
          if(counter==10'd399 )
          begin
          cir_lt_r1<=cir_lt101;
          cir_lt_r2<=cir_lt102;
          cir_lt_r3<=cir_lt103;
          cir_lt_r4<=cir_lt104;
          end
          if(counter==10'd415 )
          begin
          cir_lt_r1<=cir_lt105;
          cir_lt_r2<=cir_lt106;
          cir_lt_r3<=cir_lt107;
          cir_lt_r4<=cir_lt108;
          end
          if(counter==10'd431 )
          begin
          cir_lt_r1<=cir_lt109;
          cir_lt_r2<=cir_lt110;
          cir_lt_r3<=cir_lt111;
          cir_lt_r4<=cir_lt112;
          end
          if(counter==10'd447 )
          begin
          cir_lt_r1<=cir_lt113;
          cir_lt_r2<=cir_lt114;
          cir_lt_r3<=cir_lt115;
          cir_lt_r4<=cir_lt116;
          end
          if(counter==10'd463 )
          begin
          cir_lt_r1<=cir_lt117;
          cir_lt_r2<=cir_lt118;
          cir_lt_r3<=cir_lt119;
          cir_lt_r4<=cir_lt120;
          end
          if(counter==10'd479 )
          begin
          cir_lt_r1<=cir_lt121;
          cir_lt_r2<=cir_lt122;
          cir_lt_r3<=cir_lt123;
          cir_lt_r4<=cir_lt124;
          end
          if(counter==10'd495 )
          begin
          cir_lt_r1<=cir_lt125;
          cir_lt_r2<=cir_lt126;
          cir_lt_r3<=cir_lt127;
          cir_lt_r4<=cir_lt128;
          end
          if(counter==10'd511 )
          begin
          cir_lt_r1<=cir_lt129;
          cir_lt_r2<=cir_lt130;
          cir_lt_r3<=cir_lt131;
          cir_lt_r4<=cir_lt132;
          end
          if(counter==10'd527 )
          begin
          cir_lt_r1<=cir_lt133;
          cir_lt_r2<=cir_lt134;
          cir_lt_r3<=cir_lt135;
          cir_lt_r4<=cir_lt136;
          end
           if(counter==10'd543 )
          begin
          cir_lt_r1<=cir_lt137;
          cir_lt_r2<=cir_lt138;
          cir_lt_r3<=cir_lt139;
          cir_lt_r4<=cir_lt140;
          end
           if(counter==10'd559 )
          begin
          cir_lt_r1<=cir_lt141;
          cir_lt_r2<=cir_lt142;
          cir_lt_r3<=cir_lt143;
          cir_lt_r4<=cir_lt144;
          end
      end
    end
    dataout:
    begin
      state     <=(counter==10'd64) ? idle : dataout;
      counter   <=(counter==10'd64) ? 0    : counter+1;
      encode_fin<=1;
    end
    default:
    begin
      state     <=idle;
      counter   <=0;
      encode_fin<=1;
    end
    endcase
  end
end

endmodule

module LDPCDECg5p16v8(
                   CLK,RESET_N,start_ldpc,start_Ldata,maxiter,
                   chdata,
                   hb_count,
                   hardbit,
                   enga_en,dec_fin,dec_fail,hb_vlid,
                   ch_counta,ch_countb,addr_count);

input         CLK,RESET_N,start_ldpc,start_Ldata;
input  [4:0] maxiter;
input  [47:0] chdata;
output [3:0]  hb_count;
output [3:0]  addr_count;
output [15:0] hardbit;
output        enga_en,dec_fin,dec_fail,hb_vlid;
output [12:0] ch_counta,ch_countb;
parameter max_iter=8;
wire        data_wrsa,data_wrsb,
            deca_en,decb_en,hb_en,hb_vlid,
            load_data_en,
            memwra_en,memwrb_en,
            start_ldpc,dec_fin,vncn_en;
wire        enga_en=data_wrsa;
wire [3:0]  hb_count;
wire [3:0]  addr_count,addr_ch_count;
wire [12:0] ch_counta,ch_countb;
wire [1:0]  layer_i,section,section_r,section_ch,section_hb;
wire [4:0]  iter_count;
wire [3:0]  vncn_count;

wire [1:0] min1,min2,min3,min4,min5,min6,min7,min8,
           min9,min10,min11,min12,min13,min14,min15,min16,
           min17,min18,min19,min20,min21,min22,min23,min24,
           min25,min26,min27,min28,min29,min30,min31,min32,
           min33,min34,min35,min36,min37,min38,min39,min40,
           min41,min42,min43,min44,min45,min46,min47,min48,
           min49,min50,min51,min52,min53,min54,min55,min56,
           min57,min58,min59,min60,min61,min62,min63,min64,
           min65,min66,min67,min68,min69,min70,min71,min72,
           min73,min74,min75,min76,min77,min78,min79,min80;
wire [31:0] hbout1,hbout2,hbout3,hbout4,hbout5;
wire [15:0] hbout_o;
wire [15:0] sgn1,sgn2,sgn3,sgn4,sgn5;

wire [15:0] sgn_i=sgn1^sgn2^sgn3^sgn4^sgn5;
reg         parity_reg,dec_fail,tmn;
wire [7:0] rotat_en1,rotat_en2,rotat_en3,
           rotat_en4,rotat_en5;
reg [7:0]  rotat_en1_r,rotat_en2_r,rotat_en3_r,
           rotat_en4_r,rotat_en5_r;
always @(negedge RESET_N or posedge CLK)
begin
  if (~RESET_N)
  begin
    parity_reg<=0;
    dec_fail  <=0;
    tmn       <=0;
    rotat_en1_r <=0;
    rotat_en2_r <=0;
    rotat_en3_r <=0;
    rotat_en4_r <=0;
    rotat_en5_r <=0;
  end
  else
  begin
    tmn<= (iter_count==3'd0 & ~( vncn_count==4'd11 & addr_count==4'd15 & layer_i==2'd3))?
           1'b0 :
           (vncn_count==4'd11 & addr_count==4'd15 & layer_i==2'd3)?
           ~(parity_reg):tmn;
   if(vncn_count>4'd4)
    parity_reg<=parity_reg | sgn_i[0]
                | sgn_i[1] | sgn_i[2]
                | sgn_i[3] | sgn_i[4]
                | sgn_i[5] | sgn_i[6]
                | sgn_i[7] | sgn_i[8]
                | sgn_i[9] | sgn_i[10]
                | sgn_i[11] | sgn_i[12]
                | sgn_i[13] | sgn_i[14]
                | sgn_i[15] ;

    if(addr_count==4'd0 && layer_i==2'd0 )
      parity_reg<=0;// reset parity_reg
    if(addr_count==4'd15 && layer_i==2'd3 && iter_count==3'd7)
      dec_fail  <=parity_reg;
    rotat_en1_r <=rotat_en1;
    rotat_en2_r <=rotat_en2;
    rotat_en3_r <=rotat_en3;
    rotat_en4_r <=rotat_en4;
    rotat_en5_r <=rotat_en5;
  end
end
wire [2:0]  memgroup_hb;
wire [15:0] hardbit=hbout_o;

wire [31:0] hbout_w= (memgroup_hb==3'd0)? hbout1:
                     (memgroup_hb==3'd1)? hbout2:
                     (memgroup_hb==3'd2)? hbout3:
                     (memgroup_hb==3'd3)? hbout4: hbout5;

wire        hboutmux;
wire [15:0] hbout=(hboutmux)? hbout_w[31:16] : hbout_w[15:0];
wire [47:0] chdata, chdata_o;
wire [2:0]  memid;
wire [2:0]  memgroup;
wire [4:0] minaddrtop1,minaddrtop2,minaddrtop3,minaddrtop4,
           minaddrtop5,minaddrtop6,minaddrtop7,minaddrtop8,
           minaddrtop9,minaddrtop10,minaddrtop11,minaddrtop12,
           minaddrtop13,minaddrtop14,minaddrtop15,minaddrtop16;
wire [1:0] secmintop1,secmintop2,secmintop3,secmintop4,
           secmintop5,secmintop6,secmintop7,secmintop8,
           secmintop9,secmintop10,secmintop11,secmintop12,
           secmintop13,secmintop14,secmintop15,secmintop16,
           mintop1,mintop2,mintop3,mintop4,
           mintop5,mintop6,mintop7,mintop8,
           mintop9,mintop10,mintop11,mintop12,
           mintop13,mintop14,mintop15,mintop16;
wire [79:0] mtv1,mtv2,
            mtv9,mtv10,
            mtv17,mtv18,
            mtv25,mtv26,
            mtv33,mtv34,
            mtv1_w,mtv2_w,
            mtv9_w,mtv10_w,
            mtv17_w,mtv18_w,
            mtv25_w,mtv26_w,
            mtv33_w,mtv34_w;
wire [79:0] sumdata1,sumdata2,
            sumdata9,sumdata10,
            sumdata17,sumdata18,
            sumdata25,sumdata26,
            sumdata33,sumdata34,
            sumdata1_w,sumdata2_w,
            sumdata9_w,sumdata10_w,
            sumdata17_w,sumdata18_w,
            sumdata25_w,sumdata26_w,
            sumdata33_w,sumdata34_w;
wire [16:1]
  min_loc1 ={(minaddrtop16[0]),(minaddrtop15[0]),
             (minaddrtop14[0]),(minaddrtop13[0]),
             (minaddrtop12[0]),(minaddrtop11[0]),
             (minaddrtop10[0]),(minaddrtop9 [0]),
             (minaddrtop8 [0]),(minaddrtop7 [0]),
             (minaddrtop6 [0]),(minaddrtop5 [0]),
             (minaddrtop4 [0]),(minaddrtop3 [0]),
             (minaddrtop2 [0]),(minaddrtop1 [0])},
  min_loc2 ={(minaddrtop16[1]),(minaddrtop15[1]),
             (minaddrtop14[1]),(minaddrtop13[1]),
             (minaddrtop12[1]),(minaddrtop11[1]),
             (minaddrtop10[1]),(minaddrtop9 [1]),
             (minaddrtop8 [1]),(minaddrtop7 [1]),
             (minaddrtop6 [1]),(minaddrtop5 [1]),
             (minaddrtop4 [1]),(minaddrtop3 [1]),
             (minaddrtop2 [1]),(minaddrtop1 [1])},
  min_loc3 ={(minaddrtop16[2]),(minaddrtop15[2]),
             (minaddrtop14[2]),(minaddrtop13[2]),
             (minaddrtop12[2]),(minaddrtop11[2]),
             (minaddrtop10[2]),(minaddrtop9 [2]),
             (minaddrtop8 [2]),(minaddrtop7 [2]),
             (minaddrtop6 [2]),(minaddrtop5 [2]),
             (minaddrtop4 [2]),(minaddrtop3 [2]),
             (minaddrtop2 [2]),(minaddrtop1 [2])},
  min_loc4 ={(minaddrtop16[3]),(minaddrtop15[3]),
             (minaddrtop14[3]),(minaddrtop13[3]),
             (minaddrtop12[3]),(minaddrtop11[3]),
             (minaddrtop10[3]),(minaddrtop9 [3]),
             (minaddrtop8 [3]),(minaddrtop7 [3]),
             (minaddrtop6 [3]),(minaddrtop5 [3]),
             (minaddrtop4 [3]),(minaddrtop3 [3]),
             (minaddrtop2 [3]),(minaddrtop1 [3])},
  min_loc5 ={(minaddrtop16[4]),(minaddrtop15[4]),
             (minaddrtop14[4]),(minaddrtop13[4]),
             (minaddrtop12[4]),(minaddrtop11[4]),
             (minaddrtop10[4]),(minaddrtop9 [4]),
             (minaddrtop8 [4]),(minaddrtop7 [4]),
             (minaddrtop6 [4]),(minaddrtop5 [4]),
             (minaddrtop4 [4]),(minaddrtop3 [4]),
             (minaddrtop2 [4]),(minaddrtop1 [4])};

wire [47:0] ctm1,ctm2,ctm3,ctm4,ctm5,
            ctm6,ctm7,ctm8,ctm9,ctm10,
            ctm1_w,ctm2_w,ctm3_w,ctm4_w,
            ctm5_w,ctm6_w,ctm7_w,ctm8_w,
            ctm9_w,ctm10_w;
wire grouploaddata_en1=(memgroup==3'd0) & load_data_en,
     grouploaddata_en2=(memgroup==3'd1) & load_data_en,
     grouploaddata_en3=(memgroup==3'd2) & load_data_en,
     grouploaddata_en4=(memgroup==3'd3) & load_data_en,
     grouploaddata_en5=(memgroup==3'd4) & load_data_en;

invrotatreg invrotatreg(
                 .RESET_N(RESET_N),
                 .CLK(CLK),
                 .start_ldpc(start_ldpc),
                 .hb_en(hb_en),
                 .data_wrsa(data_wrsa),
                 .data_wrsb(data_wrsb),
                 .hbout(hbout),
                 .hbout_o(hbout_o) );

controller controller(
                     .RESET_N(RESET_N),
                     .CLK(CLK),
                     .tmn(tmn),
                     .start_ldpc(start_ldpc),
                     .maxiter(maxiter),
                     .start_Ldata(start_Ldata),
                     .data_wrsa(data_wrsa),
                     .data_wrsb(data_wrsb),
                     .deca_en(deca_en),
                     .decb_en(decb_en),
                     .hb_vlid(hb_vlid),
                     .hb_en(hb_en),
                     .load_data_en(load_data_en),
                     .dec_fin(dec_fin),
                     .vncn_en(vncn_en),
                     .memwra_en(memwra_en),
                     .memwrb_en(memwrb_en),
                     .layer_i(layer_i),
                     .section(section),
                     .section_r(section_r),
                     .iter_count(iter_count),
                     .vncn_count(vncn_count),
                     .ch_counta(ch_counta),
                     .ch_countb(ch_countb),
                     .addr_count(addr_count),
                     .addr_ch_count(addr_ch_count),
                     .hb_count(hb_count),
                     .hboutmux(hboutmux),
                     .memgroup_hb(memgroup_hb),
                     .section_hb(section_hb) );

rotatreg rotatreg(
                 .RESET_N(RESET_N),
                 .CLK(CLK),
                 .start_Ldata(start_Ldata),
                 .load_data_en(load_data_en),
                 .data_wrsa(data_wrsa),
                 .data_wrsb(data_wrsb),
                 .chdata(chdata),
                 .chdata_o(chdata_o),
                 .memid(memid),
                 .memgroup(memgroup),
                 .section_ch(section_ch) );



wire [3:0] circulant1  =4'd0 ;  //0      0       0
wire [3:0] circulant2  =4'd15;  //63      15       3
wire [3:0] circulant3  =4'd15;  //191      15       11
wire [3:0] circulant4  =4'd11;  //155      11       9
wire [3:0] circulant5  =4'd7 ;  //23      7       1
wire [3:0] circulant6  =4'd1 ;  //97      1       6
wire [3:0] circulant7  =4'd5 ;  //197      5       12
wire [3:0] circulant8  =4'd10;  //58      10       3
wire [3:0] circulant9  =4'd0 ;  //0      0       0
wire [3:0] circulant10 =4'd5 ;  //213      5       13
wire [3:0] circulant11 =4'd0 ;  //112      0       7
wire [3:0] circulant12 =4'd13;  //141      13       8
wire [3:0] circulant13 =4'd5 ;  //101      5       6
wire [3:0] circulant14 =4'd5 ;  //53      5       3
wire [3:0] circulant15 =4'd1 ;  //209      1       13
wire [3:0] circulant16 =4'd2 ;  //146      2       9
wire [3:0] circulant17 =4'd0 ;  //0      0       0
wire [3:0] circulant18 =4'd7 ;  //231      7       14
wire [3:0] circulant19 =4'd6 ;  //198      6       12
wire [3:0] circulant20 =4'd6 ;  //214      6       13
wire [3:0] circulant21 =4'd6 ;  //54      6       3
wire [3:0] circulant22 =4'd13;  //253      13       15
wire [3:0] circulant23 =4'd10;  //106      10       6
wire [3:0] circulant24 =4'd4 ;  //244      4       15

wire [3:0] circulant25 =4'd15;  //95      15       5
wire [3:0] circulant26 =4'd8 ;  //120      8       7
wire [3:0] circulant27 =4'd2 ;  //82      2       5
wire [3:0] circulant28 =4'd8 ;  //24      8       1
wire [3:0] circulant29 =4'd3 ;  //3      3       0
wire [3:0] circulant30 =4'd2 ;  //146      2       9
wire [3:0] circulant31 =4'd9 ;  //153      9       9
wire [3:0] circulant32 =4'd2 ;  //194      2       12
wire [3:0] circulant33 =4'd10;  //250      10       15
wire [3:0] circulant34 =4'd11;  //171      11       10
wire [3:0] circulant35 =4'd11;  //27      11       1
wire [3:0] circulant36 =4'd7 ;  //247      7       15
wire [3:0] circulant37 =4'd5 ;  //101      5       6
wire [3:0] circulant38 =4'd14;  //222      14       13
wire [3:0] circulant39 =4'd1 ;  //145      1       9
wire [3:0] circulant40 =4'd1 ;  //33      1       2
wire [3:0] circulant41 =4'd9 ;  //233      9       14
wire [3:0] circulant42 =4'd10;  //10      10       0
wire [3:0] circulant43 =4'd13;  //205      13       12
wire [3:0] circulant44 =4'd13;  //189      13       11
wire [3:0] circulant45 =4'd12;  //28      12       1
wire [3:0] circulant46 =4'd12;  //124      12       7
wire [3:0] circulant47 =4'd2 ;  //66      2       4
wire [3:0] circulant48 =4'd13;  //221      13       13

wire [3:0] circulant49 =4'd5 ;  //229      5       14
wire [3:0] circulant50 =4'd12;  //12      12       0
wire [3:0] circulant51 =4'd2 ;  //210      2       13
wire [3:0] circulant52 =4'd9 ;  //73      9       4
wire [3:0] circulant53 =4'd0 ;  //0      0       0
wire [3:0] circulant54 =4'd13;  //141      13       8
wire [3:0] circulant55 =4'd10;  //58      10       3
wire [3:0] circulant56 =4'd15;  //15      15       0
wire [3:0] circulant57 =4'd11;  //75      11       4
wire [3:0] circulant58 =4'd6 ;  //230      6       14
wire [3:0] circulant59 =4'd7 ;  //231      7       14
wire [3:0] circulant60 =4'd15;  //127      15       7
wire [3:0] circulant61 =4'd1 ;  //49      1       3
wire [3:0] circulant62 =4'd4 ;  //196      4       12
wire [3:0] circulant63 =4'd14;  //78      14       4
wire [3:0] circulant64 =4'd12;  //44      12       2
wire [3:0] circulant65 =4'd9 ;  //25      9       1
wire [3:0] circulant66 =4'd3 ;  //35      3       2
wire [3:0] circulant67 =4'd9 ;  //57      9       3
wire [3:0] circulant68 =4'd13;  //237      13       14
wire [3:0] circulant69 =4'd5 ;  //69      5       4
wire [3:0] circulant70 =4'd7 ;  //23      7       1
wire [3:0] circulant71 =4'd6 ;  //166      6       10
wire [3:0] circulant72 =4'd1 ;  //97      1       6

wire [3:0] circulant73 =4'd12;  //12      12       0
wire [3:0] circulant74 =4'd8 ;  //216      8       13
wire [3:0] circulant75 =4'd8 ;  //216      8       13
wire [3:0] circulant76 =4'd8 ;  //200      8       12
wire [3:0] circulant77 =4'd13;  //109      13       6
wire [3:0] circulant78 =4'd11;  //43      11       2
wire [3:0] circulant79 =4'd13;  //189      13       11
wire [3:0] circulant80 =4'd0 ;  //208      0       13
wire [3:0] circulant81 =4'd2 ;  //130      2       8
wire [3:0] circulant82 =4'd4 ;  //68      4       4
wire [3:0] circulant83 =4'd9 ;  //121      9       7
wire [3:0] circulant84 =4'd11;  //139      11       8
wire [3:0] circulant85 =4'd5 ;  //69      5       4
wire [3:0] circulant86 =4'd2 ;  //242      2       15
wire [3:0] circulant87 =4'd10;  //154      10       9
wire [3:0] circulant88 =4'd2 ;  //162      2       10
wire [3:0] circulant89 =4'd7 ;  //55      7       3
wire [3:0] circulant90 =4'd9 ;  //41      9       2
wire [3:0] circulant91 =4'd6 ;  //54      6       3
wire [3:0] circulant92 =4'd13;  //13      13       0
wire [3:0] circulant93 =4'd13;  //45      13       2
wire [3:0] circulant94 =4'd15;  //47      15       2
wire [3:0] circulant95 =4'd0 ;  //224      0       14
wire [3:0] circulant96 =4'd7 ;  //119      7       7

wire [3:0] circulant97 =4'd3 ;  //179      3       11
wire [3:0] circulant98 =4'd8 ;  //72      8       4
wire [3:0] circulant99 =4'd0 ;  //160      0       10
wire [3:0] circulant100=4'd9 ;  //89      9       5
wire [3:0] circulant101=4'd14;  //62      14       3
wire [3:0] circulant102=4'd1 ;  //49      1       3
wire [3:0] circulant103=4'd3 ;  //67      3       4
wire [3:0] circulant104=4'd5 ;  //133      5       8
wire [3:0] circulant105=4'd8 ;  //184      8       11
wire [3:0] circulant106=4'd10;  //218      10       13
wire [3:0] circulant107=4'd9 ;  //9      9       0
wire [3:0] circulant108=4'd0 ;  //80      0       5
wire [3:0] circulant109=4'd11;  //43      11       2
wire [3:0] circulant110=4'd14;  //14      14       0
wire [3:0] circulant111=4'd11;  //27      11       1
wire [3:0] circulant112=4'd10;  //170      10       10
wire [3:0] circulant113=4'd15;  //191      15       11
wire [3:0] circulant114=4'd4 ;  //228      4       14
wire [3:0] circulant115=4'd9 ;  //201      9       12
wire [3:0] circulant116=4'd6 ;  //102      6       6
wire [3:0] circulant117=4'd6 ;  //198      6       12
wire [3:0] circulant118=4'd13;  //125      13       7
wire [3:0] circulant119=4'd13;  //141      13       8
wire [3:0] circulant120=4'd4 ;  //100      4       6

wire [3:0]
  addr_count1_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant1:
                 (layer_i==2'b10)? addr_count+circulant9 :
                                   addr_count+circulant17 ,
  addr_count1_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant2:
                 (layer_i==2'b10)? addr_count+circulant10:
                                   addr_count+circulant18,
  addr_count1_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant3:
                 (layer_i==2'b10)? addr_count+circulant11:
                                   addr_count+circulant19,
  addr_count1_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant4:
                 (layer_i==2'b10)? addr_count+circulant12:
                                   addr_count+circulant20,
  addr_count2_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant5:
                 (layer_i==2'b10)? addr_count+circulant13:
                                   addr_count+circulant21,
  addr_count2_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant6:
                 (layer_i==2'b10)? addr_count+circulant14:
                                   addr_count+circulant22,
  addr_count2_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant7:
                 (layer_i==2'b10)? addr_count+circulant15:
                                   addr_count+circulant23,
  addr_count2_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant8:
                 (layer_i==2'b10)? addr_count+circulant16:
                                   addr_count+circulant24,

  addr_count3_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant25:
                 (layer_i==2'b10)? addr_count+circulant33 :
                                   addr_count+circulant41 ,
  addr_count3_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant26:
                 (layer_i==2'b10)? addr_count+circulant34:
                                   addr_count+circulant42,
  addr_count3_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant27:
                 (layer_i==2'b10)? addr_count+circulant35:
                                   addr_count+circulant43,
  addr_count3_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant28:
                 (layer_i==2'b10)? addr_count+circulant36:
                                   addr_count+circulant44,
  addr_count4_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant29:
                 (layer_i==2'b10)? addr_count+circulant37:
                                   addr_count+circulant45,
  addr_count4_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant30:
                 (layer_i==2'b10)? addr_count+circulant38:
                                   addr_count+circulant46,
  addr_count4_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant31:
                 (layer_i==2'b10)? addr_count+circulant39:
                                   addr_count+circulant47,
  addr_count4_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant32:
                 (layer_i==2'b10)? addr_count+circulant40:
                                   addr_count+circulant48,

  addr_count5_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant49:
                 (layer_i==2'b10)? addr_count+circulant57:
                                   addr_count+circulant65 ,
  addr_count5_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant50:
                 (layer_i==2'b10)? addr_count+circulant58:
                                   addr_count+circulant66,
  addr_count5_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant51:
                 (layer_i==2'b10)? addr_count+circulant59:
                                   addr_count+circulant67,
  addr_count5_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant52:
                 (layer_i==2'b10)? addr_count+circulant60:
                                   addr_count+circulant68,
  addr_count6_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant53:
                 (layer_i==2'b10)? addr_count+circulant61:
                                   addr_count+circulant69,
  addr_count6_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant54:
                 (layer_i==2'b10)? addr_count+circulant62:
                                   addr_count+circulant70,
  addr_count6_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant55:
                 (layer_i==2'b10)? addr_count+circulant63:
                                   addr_count+circulant71,
  addr_count6_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant56:
                 (layer_i==2'b10)? addr_count+circulant64:
                                   addr_count+circulant72,

  addr_count7_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant73:
                 (layer_i==2'b10)? addr_count+circulant81:
                                   addr_count+circulant89 ,
  addr_count7_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant74:
                 (layer_i==2'b10)? addr_count+circulant82:
                                   addr_count+circulant90,
  addr_count7_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant75:
                 (layer_i==2'b10)? addr_count+circulant83:
                                   addr_count+circulant91,
  addr_count7_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant76:
                 (layer_i==2'b10)? addr_count+circulant84:
                                   addr_count+circulant92,
  addr_count8_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant77:
                 (layer_i==2'b10)? addr_count+circulant85:
                                   addr_count+circulant93,
  addr_count8_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant78:
                 (layer_i==2'b10)? addr_count+circulant86:
                                   addr_count+circulant94,
  addr_count8_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant79:
                 (layer_i==2'b10)? addr_count+circulant87:
                                   addr_count+circulant95,
  addr_count8_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant80:
                 (layer_i==2'b10)? addr_count+circulant88:
                                   addr_count+circulant96,

  addr_count9_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant97:
                 (layer_i==2'b10)? addr_count+circulant105:
                                   addr_count+circulant113,
  addr_count9_2= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant98:
                 (layer_i==2'b10)? addr_count+circulant106:
                                   addr_count+circulant114,
  addr_count9_3= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant99:
                 (layer_i==2'b10)? addr_count+circulant107:
                                   addr_count+circulant115,
  addr_count9_4= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant100:
                 (layer_i==2'b10)? addr_count+circulant108:
                                   addr_count+circulant116,
  addr_count10_1= (layer_i==2'b00)? addr_count:
                 (layer_i==2'b01)? addr_count+circulant101:
                 (layer_i==2'b10)? addr_count+circulant109:
                                   addr_count+circulant117,
  addr_count10_2= (layer_i==2'b00)? addr_count:
                  (layer_i==2'b01)? addr_count+circulant102:
                  (layer_i==2'b10)? addr_count+circulant110:
                                    addr_count+circulant118,
  addr_count10_3= (layer_i==2'b00)? addr_count:
                  (layer_i==2'b01)? addr_count+circulant103:
                  (layer_i==2'b10)? addr_count+circulant111:
                                    addr_count+circulant119,
  addr_count10_4= (layer_i==2'b00)? addr_count:
                  (layer_i==2'b01)? addr_count+circulant104:
                  (layer_i==2'b10)? addr_count+circulant112:
                                    addr_count+circulant120;


assign
  rotat_en1[0]  = ((addr_count1_1  < circulant1  ) & (layer_i==2'b01)) |
                  ((addr_count1_1  < circulant9  ) & (layer_i==2'b10)) |
                  ((addr_count1_1  < circulant17 ) & (layer_i==2'b11)),
  rotat_en1[1]  = ((addr_count1_2  < circulant2  ) & (layer_i==2'b01)) |
                  ((addr_count1_2  < circulant10 ) & (layer_i==2'b10)) |
                  ((addr_count1_2  < circulant18 ) & (layer_i==2'b11)),
  rotat_en1[2]  = ((addr_count1_3  < circulant3  ) & (layer_i==2'b01)) |
                  ((addr_count1_3  < circulant11 ) & (layer_i==2'b10)) |
                  ((addr_count1_3  < circulant19 ) & (layer_i==2'b11)),
  rotat_en1[3]  = ((addr_count1_4  < circulant4  ) & (layer_i==2'b01)) |
                  ((addr_count1_4  < circulant12 ) & (layer_i==2'b10)) |
                  ((addr_count1_4  < circulant20 ) & (layer_i==2'b11)),
  rotat_en1[4]  = ((addr_count2_1  < circulant5  ) & (layer_i==2'b01)) |
                  ((addr_count2_1  < circulant13 ) & (layer_i==2'b10)) |
                  ((addr_count2_1  < circulant21 ) & (layer_i==2'b11)),
  rotat_en1[5]  = ((addr_count2_2  < circulant6  ) & (layer_i==2'b01)) |
                  ((addr_count2_2  < circulant14 ) & (layer_i==2'b10)) |
                  ((addr_count2_2  < circulant22 ) & (layer_i==2'b11)),
  rotat_en1[6]  = ((addr_count2_3  < circulant7  ) & (layer_i==2'b01)) |
                  ((addr_count2_3  < circulant15 ) & (layer_i==2'b10)) |
                  ((addr_count2_3  < circulant23 ) & (layer_i==2'b11)),
  rotat_en1[7]  = ((addr_count2_4  < circulant8  ) & (layer_i==2'b01)) |
                  ((addr_count2_4  < circulant16 ) & (layer_i==2'b10)) |
                  ((addr_count2_4  < circulant24 ) & (layer_i==2'b11)),
  rotat_en2[0]  = ((addr_count3_1  < circulant25 ) & (layer_i==2'b01)) |
                  ((addr_count3_1  < circulant33 ) & (layer_i==2'b10)) |
                  ((addr_count3_1  < circulant41 ) & (layer_i==2'b11)),
  rotat_en2[1]  = ((addr_count3_2  < circulant26 ) & (layer_i==2'b01)) |
                  ((addr_count3_2  < circulant34 ) & (layer_i==2'b10)) |
                  ((addr_count3_2  < circulant42 ) & (layer_i==2'b11)),
  rotat_en2[2]  = ((addr_count3_3  < circulant27 ) & (layer_i==2'b01)) |
                  ((addr_count3_3  < circulant35 ) & (layer_i==2'b10)) |
                  ((addr_count3_3  < circulant43 ) & (layer_i==2'b11)),
  rotat_en2[3]  = ((addr_count3_4  < circulant28 ) & (layer_i==2'b01)) |
                  ((addr_count3_4  < circulant36 ) & (layer_i==2'b10)) |
                  ((addr_count3_4  < circulant44 ) & (layer_i==2'b11)),
  rotat_en2[4]  = ((addr_count4_1  < circulant29 ) & (layer_i==2'b01)) |
                  ((addr_count4_1  < circulant37 ) & (layer_i==2'b10)) |
                  ((addr_count4_1  < circulant45 ) & (layer_i==2'b11)),
  rotat_en2[5]  = ((addr_count4_2  < circulant30 ) & (layer_i==2'b01)) |
                  ((addr_count4_2  < circulant38 ) & (layer_i==2'b10)) |
                  ((addr_count4_2  < circulant46 ) & (layer_i==2'b11)),
  rotat_en2[6]  = ((addr_count4_3  < circulant31 ) & (layer_i==2'b01)) |
                  ((addr_count4_3  < circulant39 ) & (layer_i==2'b10)) |
                  ((addr_count4_3  < circulant47 ) & (layer_i==2'b11)),
  rotat_en2[7]  = ((addr_count4_4  < circulant32 ) & (layer_i==2'b01)) |
                  ((addr_count4_4  < circulant40 ) & (layer_i==2'b10)) |
                  ((addr_count4_4  < circulant48 ) & (layer_i==2'b11)),
  rotat_en3[0]  = ((addr_count5_1  < circulant49 ) & (layer_i==2'b01)) |
                  ((addr_count5_1  < circulant57 ) & (layer_i==2'b10)) |
                  ((addr_count5_1  < circulant65 ) & (layer_i==2'b11)),
  rotat_en3[1]  = ((addr_count5_2  < circulant50 ) & (layer_i==2'b01)) |
                  ((addr_count5_2  < circulant58 ) & (layer_i==2'b10)) |
                  ((addr_count5_2  < circulant66 ) & (layer_i==2'b11)),
  rotat_en3[2]  = ((addr_count5_3  < circulant51 ) & (layer_i==2'b01)) |
                  ((addr_count5_3  < circulant59 ) & (layer_i==2'b10)) |
                  ((addr_count5_3  < circulant67 ) & (layer_i==2'b11)),
  rotat_en3[3]  = ((addr_count5_4  < circulant52 ) & (layer_i==2'b01)) |
                  ((addr_count5_4  < circulant60 ) & (layer_i==2'b10)) |
                  ((addr_count5_4  < circulant68 ) & (layer_i==2'b11)),
  rotat_en3[4]  = ((addr_count6_1  < circulant53 ) & (layer_i==2'b01)) |
                  ((addr_count6_1  < circulant61 ) & (layer_i==2'b10)) |
                  ((addr_count6_1  < circulant69 ) & (layer_i==2'b11)),
  rotat_en3[5]  = ((addr_count6_2  < circulant54 ) & (layer_i==2'b01)) |
                  ((addr_count6_2  < circulant62 ) & (layer_i==2'b10)) |
                  ((addr_count6_2  < circulant70 ) & (layer_i==2'b11)),
  rotat_en3[6]  = ((addr_count6_3  < circulant55 ) & (layer_i==2'b01)) |
                  ((addr_count6_3  < circulant63 ) & (layer_i==2'b10)) |
                  ((addr_count6_3  < circulant71 ) & (layer_i==2'b11)),
  rotat_en3[7]  = ((addr_count6_4  < circulant56 ) & (layer_i==2'b01)) |
                  ((addr_count6_4  < circulant64 ) & (layer_i==2'b10)) |
                  ((addr_count6_4  < circulant72 ) & (layer_i==2'b11)),
  rotat_en4[0]  = ((addr_count7_1  < circulant73 ) & (layer_i==2'b01)) |
                  ((addr_count7_1  < circulant81 ) & (layer_i==2'b10)) |
                  ((addr_count7_1  < circulant89 ) & (layer_i==2'b11)),
  rotat_en4[1]  = ((addr_count7_2  < circulant74 ) & (layer_i==2'b01)) |
                  ((addr_count7_2  < circulant82 ) & (layer_i==2'b10)) |
                  ((addr_count7_2  < circulant90 ) & (layer_i==2'b11)),
  rotat_en4[2]  = ((addr_count7_3  < circulant75 ) & (layer_i==2'b01)) |
                  ((addr_count7_3  < circulant83 ) & (layer_i==2'b10)) |
                  ((addr_count7_3  < circulant91 ) & (layer_i==2'b11)),
  rotat_en4[3]  = ((addr_count7_4  < circulant76 ) & (layer_i==2'b01)) |
                  ((addr_count7_4  < circulant84 ) & (layer_i==2'b10)) |
                  ((addr_count7_4  < circulant92 ) & (layer_i==2'b11)),
  rotat_en4[4]  = ((addr_count8_1  < circulant77 ) & (layer_i==2'b01)) |
                  ((addr_count8_1  < circulant85 ) & (layer_i==2'b10)) |
                  ((addr_count8_1  < circulant93 ) & (layer_i==2'b11)),
  rotat_en4[5]  = ((addr_count8_2  < circulant78 ) & (layer_i==2'b01)) |
                  ((addr_count8_2  < circulant86 ) & (layer_i==2'b10)) |
                  ((addr_count8_2  < circulant94 ) & (layer_i==2'b11)),
  rotat_en4[6]  = ((addr_count8_3  < circulant79 ) & (layer_i==2'b01)) |
                  ((addr_count8_3  < circulant87 ) & (layer_i==2'b10)) |
                  ((addr_count8_3  < circulant95 ) & (layer_i==2'b11)),
  rotat_en4[7]  = ((addr_count8_4  < circulant80 ) & (layer_i==2'b01)) |
                  ((addr_count8_4  < circulant88 ) & (layer_i==2'b10)) |
                  ((addr_count8_4  < circulant96 ) & (layer_i==2'b11)),
  rotat_en5[0] =  ((addr_count9_1  < circulant97 ) & (layer_i==2'b01)) |
                  ((addr_count9_1  < circulant105) & (layer_i==2'b10)) |
                  ((addr_count9_1  < circulant113) & (layer_i==2'b11)),
  rotat_en5[1] =  ((addr_count9_2  < circulant98 ) & (layer_i==2'b01)) |
                  ((addr_count9_2  < circulant106) & (layer_i==2'b10)) |
                  ((addr_count9_2  < circulant114) & (layer_i==2'b11)),
  rotat_en5[2] =  ((addr_count9_3  < circulant99 ) & (layer_i==2'b01)) |
                  ((addr_count9_3  < circulant107) & (layer_i==2'b10)) |
                  ((addr_count9_3  < circulant115) & (layer_i==2'b11)),
  rotat_en5[3] =  ((addr_count9_4  < circulant100) & (layer_i==2'b01)) |
                  ((addr_count9_4  < circulant108) & (layer_i==2'b10)) |
                  ((addr_count9_4  < circulant116) & (layer_i==2'b11)),
  rotat_en5[4] =  ((addr_count10_1 < circulant101) & (layer_i==2'b01)) |
                  ((addr_count10_1 < circulant109) & (layer_i==2'b10)) |
                  ((addr_count10_1 < circulant117) & (layer_i==2'b11)),
  rotat_en5[5] =  ((addr_count10_2 < circulant102) & (layer_i==2'b01)) |
                  ((addr_count10_2 < circulant110) & (layer_i==2'b10)) |
                  ((addr_count10_2 < circulant118) & (layer_i==2'b11)),
  rotat_en5[6] =  ((addr_count10_3 < circulant103) & (layer_i==2'b01)) |
                  ((addr_count10_3 < circulant111) & (layer_i==2'b10)) |
                  ((addr_count10_3 < circulant119) & (layer_i==2'b11)),
  rotat_en5[7] =  ((addr_count10_4 < circulant104) & (layer_i==2'b01)) |
                  ((addr_count10_4 < circulant112) & (layer_i==2'b10)) |
                  ((addr_count10_4 < circulant120) & (layer_i==2'b11));

vncngroup vncngroup1(
          .CLK(CLK),.RESET_N(RESET_N),
          .start_ldpc(start_ldpc),.vncn_en(vncn_en),
          .chdata(chdata_o),
          .layer_i(layer_i),
          .section(section),.section_r(section_r),.section_ch(section_ch),.section_hb(section_hb),
          .iter_count(iter_count),
          .vncn_count(vncn_count),
          .tmn(tmn),
          .data_wrsa(data_wrsa),.data_wrsb(data_wrsb),
          .deca_en(deca_en),.decb_en(decb_en),
          .memwra_en(memwra_en),.memwrb_en(memwrb_en),
          .grouploaddata_en(grouploaddata_en1),
          .hb_count(hb_count),
          .addr_count(addr_count),.addr_ch_count(addr_ch_count),
          .memid(memid),
          .min_loc (min_loc1 ),
          .min_i1(mintop1),.min_i2(mintop2),
          .min_i3(mintop3),.min_i4(mintop4),
          .min_i5(mintop5),.min_i6(mintop6),
          .min_i7(mintop7),.min_i8(mintop8),
          .min_i9(mintop9),.min_i10(mintop10),
          .min_i11(mintop11),.min_i12(mintop12),
          .min_i13(mintop13),.min_i14(mintop14),
          .min_i15(mintop15),.min_i16(mintop16),
          .secmin_i1(secmintop1),.secmin_i2(secmintop2),
          .secmin_i3(secmintop3),.secmin_i4(secmintop4),
          .secmin_i5(secmintop5),.secmin_i6(secmintop6),
          .secmin_i7(secmintop7),.secmin_i8(secmintop8),
          .secmin_i9(secmintop9),.secmin_i10(secmintop10),
          .secmin_i11(secmintop11),.secmin_i12(secmintop12),
          .secmin_i13(secmintop13),.secmin_i14(secmintop14),
          .secmin_i15(secmintop15),.secmin_i16(secmintop16),
          .mtv1_i (mtv1_w ),.mtv2_i (mtv2_w ),
          .sumdata1_i(sumdata1_w),.sumdata2_i(sumdata2_w),                                                                               
          .ctm1_i(ctm1),.ctm2_i(ctm2),
          .addr_count1_1(addr_count1_1),.addr_count1_2(addr_count1_2),
          .addr_count1_3(addr_count1_3),.addr_count1_4(addr_count1_4),
          .addr_count2_1(addr_count2_1),.addr_count2_2(addr_count2_2),
          .addr_count2_3(addr_count2_3),.addr_count2_4(addr_count2_4),
          .hbout(hbout1),
          .min1(min1),.min2(min2),.min3(min3),.min4(min4),
          .min5(min5),.min6(min6),.min7(min7),.min8(min8),
          .min9(min9),.min10(min10),.min11(min11),.min12(min12),
          .min13(min13),.min14(min14),.min15(min15),.min16(min16),
          .sgn(sgn1),.sgn_i(sgn_i),
          .mtv1_o (mtv1 ),.mtv2_o (mtv2 ),
          .ctm1(ctm1_w),.ctm2(ctm2_w),
          .sumdata1(sumdata1),.sumdata2(sumdata2));                                                                                      


invpermutator1 invpermutator1(
               .layer_i(layer_i),.section(section_r),
               .mtv1 (mtv1 ),.mtv2 (mtv2 ),
               .mtv1_w (mtv1_w ),.mtv2_w (mtv2_w ),
               .ctm1_i(ctm1_w),.ctm2_i(ctm2_w),
               .sumdata1(sumdata1),.sumdata2(sumdata2),
               .sumdata1_w(sumdata1_w),.sumdata2_w(sumdata2_w),
               .rotat_en(rotat_en1_r),
               .ctm1(ctm1),.ctm2(ctm2) );
vncngroup vncngroup2(
          .CLK(CLK),.RESET_N(RESET_N),
          .start_ldpc(start_ldpc),.vncn_en(vncn_en),
          .chdata(chdata_o),
          .layer_i(layer_i),
          .section(section),.section_r(section_r),.section_ch(section_ch),.section_hb(section_hb),
          .iter_count(iter_count),
          .vncn_count(vncn_count),
          .tmn(tmn),
          .data_wrsa(data_wrsa),.data_wrsb(data_wrsb),
          .deca_en(deca_en),.decb_en(decb_en),
          .memwra_en(memwra_en),.memwrb_en(memwrb_en),
          .grouploaddata_en(grouploaddata_en2),
          .hb_count(hb_count),
          .addr_count(addr_count),.addr_ch_count(addr_ch_count),
          .memid(memid),
          .min_loc (min_loc2),
          .min_i1(mintop1),.min_i2(mintop2),
          .min_i3(mintop3),.min_i4(mintop4),
          .min_i5(mintop5),.min_i6(mintop6),
          .min_i7(mintop7),.min_i8(mintop8),
          .min_i9(mintop9),.min_i10(mintop10),
          .min_i11(mintop11),.min_i12(mintop12),
          .min_i13(mintop13),.min_i14(mintop14),
          .min_i15(mintop15),.min_i16(mintop16),
          .secmin_i1(secmintop1),.secmin_i2(secmintop2),
          .secmin_i3(secmintop3),.secmin_i4(secmintop4),
          .secmin_i5(secmintop5),.secmin_i6(secmintop6),
          .secmin_i7(secmintop7),.secmin_i8(secmintop8),
          .secmin_i9(secmintop9),.secmin_i10(secmintop10),
          .secmin_i11(secmintop11),.secmin_i12(secmintop12),
          .secmin_i13(secmintop13),.secmin_i14(secmintop14),
          .secmin_i15(secmintop15),.secmin_i16(secmintop16),
          .mtv1_i (mtv9_w ),.mtv2_i(mtv10_w),
          .sumdata1_i(sumdata9_w),.sumdata2_i(sumdata10_w),                                                                              
          .ctm1_i(ctm3),.ctm2_i(ctm4),
          .addr_count1_1(addr_count3_1),.addr_count1_2(addr_count3_2),
          .addr_count1_3(addr_count3_3),.addr_count1_4(addr_count3_4),
          .addr_count2_1(addr_count4_1),.addr_count2_2(addr_count4_2),
          .addr_count2_3(addr_count4_3),.addr_count2_4(addr_count4_4),
          .hbout(hbout2),
          .min1 (min17),.min2 (min18),.min3 (min19),.min4 (min20),
          .min5 (min21),.min6 (min22),.min7 (min23),.min8 (min24),
          .min9 (min25),.min10(min26),.min11(min27),.min12(min28),
          .min13(min29),.min14(min30),.min15(min31),.min16(min32),
          .sgn(sgn2),.sgn_i(sgn_i),
          .mtv1_o (mtv9 ),.mtv2_o(mtv10),
          .ctm1(ctm3_w),.ctm2(ctm4_w),
          .sumdata1(sumdata9),.sumdata2(sumdata10));                                                                                     


invpermutator2 invpermutator2(
                     .layer_i(layer_i),.section(section_r),
                     .mtv1 (mtv9 ),.mtv2(mtv10),
                     .mtv1_w (mtv9_w ),.mtv2_w(mtv10_w),
                     .ctm1_i(ctm3_w),.ctm2_i(ctm4_w),
                     .sumdata1(sumdata9),.sumdata2(sumdata10),
                     .sumdata1_w(sumdata9_w),.sumdata2_w(sumdata10_w),
                     .rotat_en(rotat_en2_r),
                     .ctm1(ctm3),.ctm2(ctm4)  );

vncngroup vncngroup3(
             .CLK(CLK),.RESET_N(RESET_N),
             .start_ldpc(start_ldpc),.vncn_en(vncn_en),
             .chdata(chdata_o),
             .layer_i(layer_i),
             .section(section),.section_r(section_r),.section_ch(section_ch),.section_hb(section_hb),
             .iter_count(iter_count),
             .vncn_count(vncn_count),
             .tmn(tmn),
             .data_wrsa(data_wrsa),.data_wrsb(data_wrsb),
             .deca_en(deca_en),.decb_en(decb_en),
             .memwra_en(memwra_en),.memwrb_en(memwrb_en),
             .grouploaddata_en(grouploaddata_en3),
             .hb_count(hb_count),
             .addr_count(addr_count),.addr_ch_count(addr_ch_count),
             .memid(memid),
             .min_loc (min_loc3 ),
             .min_i1(mintop1),.min_i2(mintop2),
             .min_i3(mintop3),.min_i4(mintop4),
             .min_i5(mintop5),.min_i6(mintop6),
             .min_i7(mintop7),.min_i8(mintop8),
             .min_i9(mintop9),.min_i10(mintop10),
             .min_i11(mintop11),.min_i12(mintop12),
             .min_i13(mintop13),.min_i14(mintop14),
             .min_i15(mintop15),.min_i16(mintop16),
             .secmin_i1(secmintop1),.secmin_i2(secmintop2),
             .secmin_i3(secmintop3),.secmin_i4(secmintop4),
             .secmin_i5(secmintop5),.secmin_i6(secmintop6),
             .secmin_i7(secmintop7),.secmin_i8(secmintop8),
             .secmin_i9(secmintop9),.secmin_i10(secmintop10),
             .secmin_i11(secmintop11),.secmin_i12(secmintop12),
             .secmin_i13(secmintop13),.secmin_i14(secmintop14),
             .secmin_i15(secmintop15),.secmin_i16(secmintop16),
             .mtv1_i (mtv17_w),.mtv2_i(mtv18_w),
             .sumdata1_i(sumdata17_w),.sumdata2_i(sumdata18_w),
             .ctm1_i(ctm5),.ctm2_i(ctm6),
             .addr_count1_1(addr_count5_1),.addr_count1_2(addr_count5_2),
             .addr_count1_3(addr_count5_3),.addr_count1_4(addr_count5_4),
             .addr_count2_1(addr_count6_1),.addr_count2_2(addr_count6_2),
             .addr_count2_3(addr_count6_3),.addr_count2_4(addr_count6_4),
             .hbout(hbout3),
             .min1 (min33),.min2 (min34),.min3 (min35),.min4 (min36),
             .min5 (min37),.min6 (min38),.min7 (min39),.min8 (min40),
             .min9 (min41),.min10(min42),.min11(min43),.min12(min44),
             .min13(min45),.min14(min46),.min15(min47),.min16(min48),
             .sgn(sgn3),.sgn_i(sgn_i),
             .mtv1_o (mtv17 ),.mtv2_o (mtv18 ),
             .ctm1(ctm5_w),.ctm2(ctm6_w),
             .sumdata1(sumdata17),.sumdata2(sumdata18) );                                                                                
invpermutator3 invpermutator3(
                      .layer_i(layer_i),.section(section_r),
                      .mtv1 (mtv17 ),.mtv2 (mtv18 ),
                      .mtv1_w (mtv17_w ),.mtv2_w (mtv18_w ),
                      .ctm1_i(ctm5_w),.ctm2_i(ctm6_w),
                      .sumdata1(sumdata17),.sumdata2(sumdata18),
                      .sumdata1_w(sumdata17_w),.sumdata2_w(sumdata18_w),
                      .rotat_en(rotat_en3_r),
                      .ctm1(ctm5),.ctm2(ctm6)   );

vncngroup vncngroup4(
             .CLK(CLK),.RESET_N(RESET_N),.start_ldpc(start_ldpc),.vncn_en(vncn_en),
             .chdata(chdata_o),
             .layer_i(layer_i),
             .section(section),.section_r(section_r),.section_ch(section_ch),.section_hb(section_hb),
             .iter_count(iter_count),
             .vncn_count(vncn_count),
             .tmn(tmn),
             .data_wrsa(data_wrsa),.data_wrsb(data_wrsb),
             .deca_en(deca_en),.decb_en(decb_en),
             .memwra_en(memwra_en),.memwrb_en(memwrb_en),
             .grouploaddata_en(grouploaddata_en4),
             .hb_count(hb_count),
             .addr_count(addr_count),.addr_ch_count(addr_ch_count),
             .memid(memid),
             .min_loc (min_loc4 ),
             .min_i1(mintop1),.min_i2(mintop2),
             .min_i3(mintop3),.min_i4(mintop4),
             .min_i5(mintop5),.min_i6(mintop6),
             .min_i7(mintop7),.min_i8(mintop8),
             .min_i9(mintop9),.min_i10(mintop10),
             .min_i11(mintop11),.min_i12(mintop12),
             .min_i13(mintop13),.min_i14(mintop14),
             .min_i15(mintop15),.min_i16(mintop16),
             .secmin_i1(secmintop1),.secmin_i2(secmintop2),
             .secmin_i3(secmintop3),.secmin_i4(secmintop4),
             .secmin_i5(secmintop5),.secmin_i6(secmintop6),
             .secmin_i7(secmintop7),.secmin_i8(secmintop8),
             .secmin_i9(secmintop9),.secmin_i10(secmintop10),
             .secmin_i11(secmintop11),.secmin_i12(secmintop12),
             .secmin_i13(secmintop13),.secmin_i14(secmintop14),
             .secmin_i15(secmintop15),.secmin_i16(secmintop16),
             .mtv1_i (mtv25_w ),.mtv2_i (mtv26_w ),
             .sumdata1_i(sumdata25_w),.sumdata2_i(sumdata26_w),
             .ctm1_i(ctm7),.ctm2_i(ctm8),
             .addr_count1_1(addr_count7_1),.addr_count1_2(addr_count7_2),
             .addr_count1_3(addr_count7_3),.addr_count1_4(addr_count7_4),
             .addr_count2_1(addr_count8_1),.addr_count2_2(addr_count8_2),
             .addr_count2_3(addr_count8_3),.addr_count2_4(addr_count8_4),
             .hbout(hbout4),
             .min1 (min49),.min2 (min50),.min3 (min51),.min4 (min52),
             .min5 (min53),.min6 (min54),.min7 (min55),.min8 (min56),
             .min9 (min57),.min10(min58),.min11(min59),.min12(min60),
             .min13(min61),.min14(min62),.min15(min63),.min16(min64),
             .sgn(sgn4),.sgn_i(sgn_i),
             .mtv1_o (mtv25 ),.mtv2_o (mtv26 ),
             .ctm1(ctm7_w),.ctm2(ctm8_w),
             .sumdata1(sumdata25),.sumdata2(sumdata26) );                                                                                
invpermutator4 invpermutator4(
                      .layer_i(layer_i),.section(section_r),
                      .mtv1 (mtv25 ),.mtv2 (mtv26 ),
                      .mtv1_w (mtv25_w ),.mtv2_w (mtv26_w ),
                      .ctm1_i(ctm7_w),.ctm2_i(ctm8_w),
                      .sumdata1(sumdata25),.sumdata2(sumdata26),
                      .sumdata1_w(sumdata25_w),.sumdata2_w(sumdata26_w),
                      .rotat_en(rotat_en4_r),
                      .ctm1(ctm7),.ctm2(ctm8)  );

vncngroup vncngroup5(
             .CLK(CLK),.RESET_N(RESET_N),
             .start_ldpc(start_ldpc),.vncn_en(vncn_en),
             .chdata(chdata_o),
             .layer_i(layer_i),
             .section(section),.section_r(section_r),.section_ch(section_ch),.section_hb(section_hb),
             .iter_count(iter_count),
             .vncn_count(vncn_count),
             .tmn(tmn),
             .data_wrsa(data_wrsa),.data_wrsb(data_wrsb),
             .deca_en(deca_en),.decb_en(decb_en),
             .memwra_en(memwra_en),.memwrb_en(memwrb_en),
             .grouploaddata_en(grouploaddata_en5),
             .hb_count(hb_count),
             .addr_count(addr_count),.addr_ch_count(addr_ch_count),
             .memid(memid),
             .min_loc (min_loc5 ),
             .min_i1(mintop1),.min_i2(mintop2),
             .min_i3(mintop3),.min_i4(mintop4),
             .min_i5(mintop5),.min_i6(mintop6),
             .min_i7(mintop7),.min_i8(mintop8),
             .min_i9(mintop9),.min_i10(mintop10),
             .min_i11(mintop11),.min_i12(mintop12),
             .min_i13(mintop13),.min_i14(mintop14),
             .min_i15(mintop15),.min_i16(mintop16),
             .secmin_i1(secmintop1),.secmin_i2(secmintop2),
             .secmin_i3(secmintop3),.secmin_i4(secmintop4),
             .secmin_i5(secmintop5),.secmin_i6(secmintop6),
             .secmin_i7(secmintop7),.secmin_i8(secmintop8),
             .secmin_i9(secmintop9),.secmin_i10(secmintop10),
             .secmin_i11(secmintop11),.secmin_i12(secmintop12),
             .secmin_i13(secmintop13),.secmin_i14(secmintop14),
             .secmin_i15(secmintop15),.secmin_i16(secmintop16),
             .mtv1_i (mtv33_w ),.mtv2_i (mtv34_w ),
             .sumdata1_i(sumdata33_w),.sumdata2_i(sumdata34_w),
             .ctm1_i(ctm9),.ctm2_i(ctm10),
             .addr_count1_1(addr_count9_1),.addr_count1_2(addr_count9_2),
             .addr_count1_3(addr_count9_3),.addr_count1_4(addr_count9_4),
             .addr_count2_1(addr_count10_1),.addr_count2_2(addr_count10_2),
             .addr_count2_3(addr_count10_3),.addr_count2_4(addr_count10_4),
             .hbout(hbout5),
             .min1 (min65),.min2 (min66),.min3 (min67),.min4 (min68),
             .min5 (min69),.min6 (min70),.min7 (min71),.min8 (min72),
             .min9 (min73),.min10(min74),.min11(min75),.min12(min76),
             .min13(min77),.min14(min78),.min15(min79),.min16(min80),
             .sgn(sgn5),.sgn_i(sgn_i),
             .mtv1_o (mtv33 ),.mtv2_o (mtv34 ),
             .ctm1(ctm9_w),.ctm2(ctm10_w),
             .sumdata1(sumdata33),.sumdata2(sumdata34) );                                                                                


invpermutator5 invpermutator5(
                      .layer_i(layer_i),.section(section_r),
                      .mtv1 (mtv33 ),.mtv2 (mtv34 ),
                      .mtv1_w (mtv33_w ),.mtv2_w (mtv34_w ) ,
                      .ctm1_i(ctm9_w),.ctm2_i(ctm10_w),
                      .sumdata1(sumdata33),.sumdata2(sumdata34),
                      .sumdata1_w(sumdata33_w),.sumdata2_w(sumdata34_w),
                      .rotat_en(rotat_en5_r),
                      .ctm1(ctm9),.ctm2(ctm10) );

CMPtop CMPtop1(
   .vtc_1(min1 ), .vtc_2(min17), .vtc_3(min33),
   .vtc_4(min49), .vtc_5(min65),
   .min(mintop1),
   .secmin(secmintop1),
   .minaddr(minaddrtop1)
   );

CMPtop CMPtop2(
   .vtc_1(min2 ),.vtc_2(min18),.vtc_3(min34),
   .vtc_4(min50), .vtc_5(min66),
   .min(mintop2),
   .secmin(secmintop2),
   .minaddr(minaddrtop2)
   );
CMPtop CMPtop3(
   .vtc_1(min3 ), .vtc_2(min19), .vtc_3(min35),
   .vtc_4(min51), .vtc_5(min67),
   .min(mintop3),
   .secmin(secmintop3),
   .minaddr(minaddrtop3)
   );
CMPtop CMPtop4(
   .vtc_1(min4 ), .vtc_2(min20), .vtc_3(min36),
   .vtc_4(min52), .vtc_5(min68),
   .min(mintop4),
   .secmin(secmintop4),
   .minaddr(minaddrtop4)
   );
CMPtop CMPtop5(
   .vtc_1(min5 ), .vtc_2(min21), .vtc_3(min37),
   .vtc_4(min53), .vtc_5(min69),
   .min(mintop5),
   .secmin(secmintop5),
   .minaddr(minaddrtop5)
   );
CMPtop CMPtop6(
   .vtc_1(min6 ),.vtc_2(min22),.vtc_3(min38),
   .vtc_4(min54),.vtc_5(min70),
   .min(mintop6),
   .secmin(secmintop6),
   .minaddr(minaddrtop6)
   );
CMPtop CMPtop7(
   .vtc_1(min7 ),.vtc_2(min23),.vtc_3(min39),
   .vtc_4(min55),.vtc_5(min71),
   . min(mintop7),
   . secmin(secmintop7),
   . minaddr(minaddrtop7)
   );
CMPtop CMPtop8(
   .vtc_1(min8 ),.vtc_2(min24),.vtc_3(min40),
   .vtc_4(min56),.vtc_5(min72),
   .min(mintop8),
   .secmin(secmintop8),
   .minaddr(minaddrtop8)
   );
CMPtop CMPtop9(
   .vtc_1(min9 ),.vtc_2(min25),.vtc_3(min41),
   .vtc_4(min57),.vtc_5(min73),
   .min(mintop9),
   .secmin(secmintop9),
   .minaddr(minaddrtop9)
   );
CMPtop CMPtop10(
   .vtc_1(min10),.vtc_2(min26),.vtc_3(min42),
   .vtc_4(min58),.vtc_5(min74),
   .min(mintop10),
   .secmin(secmintop10),
   .minaddr(minaddrtop10)
   );
CMPtop CMPtop11(
   .vtc_1(min11),.vtc_2(min27),.vtc_3(min43),
   .vtc_4(min59),.vtc_5(min75),
   .min(mintop11),
   .secmin(secmintop11),
   .minaddr(minaddrtop11)
   );
CMPtop CMPtop12(
   .vtc_1(min12),.vtc_2(min28),.vtc_3(min44),
   .vtc_4(min60),.vtc_5(min76),
   .min(mintop12),
   .secmin(secmintop12),
   .minaddr(minaddrtop12)
   );
CMPtop CMPtop13(
   .vtc_1(min13),.vtc_2(min29), .vtc_3(min45),
   .vtc_4(min61), .vtc_5(min77),
   .min(mintop13),
   .secmin(secmintop13),
   .minaddr(minaddrtop13)
   );
CMPtop CMPtop14(
   .vtc_1(min14), .vtc_2(min30), .vtc_3(min46),
   .vtc_4(min62), .vtc_5(min78),
   .min(mintop14),
   .secmin(secmintop14),
   .minaddr(minaddrtop14)
   );
CMPtop CMPtop15(
   .vtc_1(min15), .vtc_2(min31), .vtc_3(min47),
   .vtc_4(min63), .vtc_5(min79),
   .min(mintop15),
   .secmin(secmintop15),
   .minaddr(minaddrtop15)
   );
CMPtop CMPtop16(
   .vtc_1(min16), .vtc_2(min32), .vtc_3(min48),
   .vtc_4(min64), .vtc_5(min80),
   .min(mintop16),
   .secmin(secmintop16),
   .minaddr(minaddrtop16)
   );
endmodule
module vncngroup(
               CLK,RESET_N,start_ldpc,vncn_en,
               chdata,
               layer_i,section,section_r,section_ch,section_hb,
               iter_count,
               vncn_count,
               tmn,
               data_wrsa,data_wrsb,
               deca_en,decb_en,
               memwra_en,memwrb_en,
               grouploaddata_en,
               hb_count,
               addr_count,addr_ch_count,
               memid,
               min_loc,
               min_i1,min_i2,min_i3,min_i4,
               min_i5,min_i6,min_i7,min_i8,
               min_i9,min_i10,min_i11,min_i12,
               min_i13,min_i14,min_i15,min_i16,
               secmin_i1,secmin_i2,secmin_i3,secmin_i4,
               secmin_i5,secmin_i6,secmin_i7,secmin_i8,
               secmin_i9,secmin_i10,secmin_i11,secmin_i12,
               secmin_i13,secmin_i14,secmin_i15,secmin_i16,
               sgn_i,
               mtv1_i,mtv2_i,
               ctm1_i,ctm2_i,
               sumdata1_i,sumdata2_i,
               addr_count1_1,addr_count1_2,
               addr_count1_3,addr_count1_4,
               addr_count2_1,addr_count2_2,
               addr_count2_3,addr_count2_4,
               hbout,
               min1,min2,min3,min4,
               min5,min6,min7,min8,
               min9,min10,min11,min12,
               min13,min14,min15,min16,sgn,
               mtv1_o,mtv2_o,
               ctm1,ctm2,
               sumdata1,sumdata2);

input        CLK,RESET_N,start_ldpc,vncn_en;
input [47:0] chdata;
input [1:0] layer_i,section,section_r,section_ch,section_hb;
input [4:0] iter_count;
input [3:0] vncn_count;
input       tmn;
input       data_wrsa,data_wrsb,deca_en,decb_en,
            memwra_en,memwrb_en,grouploaddata_en;
input [3:0] hb_count;
input [3:0] addr_count,addr_ch_count;
input [2:0] memid;
input [16:1]min_loc;
input [1:0] min_i1,min_i2,min_i3,min_i4,
            min_i5,min_i6,min_i7,min_i8,
            min_i9,min_i10,min_i11,min_i12,
            min_i13,min_i14,min_i15,min_i16,
            secmin_i1,secmin_i2,secmin_i3,secmin_i4,
            secmin_i5,secmin_i6,secmin_i7,secmin_i8,
            secmin_i9,secmin_i10,secmin_i11,secmin_i12,
            secmin_i13,secmin_i14,secmin_i15,secmin_i16;
input [16:1] sgn_i;
input [79:0] mtv1_i,mtv2_i;
input [79:0] sumdata1_i,sumdata2_i;
input [47:0] ctm1_i,ctm2_i;
input [3:0] addr_count1_1,addr_count1_2,
            addr_count1_3,addr_count1_4,
            addr_count2_1,addr_count2_2,
            addr_count2_3,addr_count2_4;
output [31:0] hbout;

output [1:0] min1,min2,min3,min4,
             min5,min6,min7,min8,
             min9,min10,min11,min12,
             min13,min14,min15,min16;
output [16:1]sgn;
output [79:0] mtv1_o,mtv2_o;
output [47:0] ctm1,ctm2;
output [79:0] sumdata1,sumdata2;
wire [1:0] min1,min2,min3,min4,
           min5,min6,min7,min8,
           min9,min10,min11,min12,
           min13,min14,min15,min16;
wire [7:0] addr1a_w, addr2a_w;
wire [2:0] ctm1_1,ctm2_1,ctm1_2,ctm2_2,
           ctm1_3,ctm2_3,ctm1_4,ctm2_4,
           ctm1_5,ctm2_5,ctm1_6,ctm2_6,
           ctm1_7,ctm2_7,ctm1_8,ctm2_8,
           ctm1_9,ctm2_9,ctm1_10,ctm2_10,
           ctm1_11,ctm2_11,ctm1_12,ctm2_12,
           ctm1_13,ctm2_13,ctm1_14,ctm2_14,
           ctm1_15,ctm2_15,ctm1_16,ctm2_16;

wire [47:0] mtv1,mtv2;

wire [79:0] sumdata1a_o,sumdata2a_o,sumdata1b_o,sumdata2b_o;

wire [31:0] sr_hb;

wire hbwra_en= memwra_en & ~tmn & (layer_i==2'd0) & deca_en;
wire hbwrb_en= memwrb_en & ~tmn & (layer_i==2'd0) & decb_en;
wire dec_en= ( deca_en | decb_en ) & ~tmn ;

wire [5:0] hb_count_w={section_hb,hb_count};
wire [5:0] hb_count_wr_w={section,addr_count};
wire [5:0] hb_counta=deca_en?hb_count_wr_w:hb_count_w;
wire [5:0] hb_countb=decb_en?hb_count_wr_w:hb_count_w;

wire [31:0] hbouta,hboutb;
wire [31:0] hbout= decb_en ? hbouta : hboutb;

memblock64x32 memh_a(
          .A(hb_counta),
         .CEN(dec_en),
         .CLK(CLK),
         .D(sr_hb),
         .WEN(hbwra_en),
         .Q(hbouta)
         );
memblock64x32 memh_b(
        .A(hb_countb),
         .CEN(dec_en),
         .CLK(CLK),
         .D(sr_hb),
         .WEN(hbwrb_en),
         .Q(hboutb)
         );
wire
  chmemwra1_en =data_wrsa?
                (memid==3'd0 | memid==3'd1 |
                 memid==3'd2 | memid==3'd3  )& grouploaddata_en:memwra_en,
  chmemwra2_en =data_wrsa?
                (memid==3'd4 | memid==3'd5 |
                 memid==3'd6 | memid==3'd7  )& grouploaddata_en:memwra_en,

  chmemwrb1_en =data_wrsb?
                (memid==3'd0 | memid==3'd1 |
                 memid==3'd2 | memid==3'd3  )& grouploaddata_en:memwrb_en,
  chmemwrb2_en =data_wrsb?
                (memid==3'd4 | memid==3'd5 |
                 memid==3'd6 | memid==3'd7  )& grouploaddata_en:memwrb_en;

wire mema_en=(dec_en | data_wrsa) & ~tmn;
wire memb_en=(dec_en | data_wrsb) & ~tmn;

wire [5:0]
  addrcha1_w =(data_wrsa)?{section_ch,addr_ch_count}:addr1a_w[5:0],
  addrcha2_w =(data_wrsa)?{section_ch,addr_ch_count}:addr2a_w[5:0],
  addrchb1_w =(data_wrsb)?{section_ch,addr_ch_count}:addr1a_w[5:0],
  addrchb2_w =(data_wrsb)?{section_ch,addr_ch_count}:addr2a_w[5:0];

wire [79:0] chdata_w={chdata[47],chdata[47],chdata[47:45],chdata[44],chdata[44],chdata[44:42],
                      chdata[41],chdata[41],chdata[41:39],chdata[38],chdata[38],chdata[38:36],
                      chdata[35],chdata[35],chdata[35:33],chdata[32],chdata[32],chdata[32:30],
                      chdata[29],chdata[29],chdata[29:27],chdata[26],chdata[26],chdata[26:24],
                      chdata[23],chdata[23],chdata[23:21],chdata[20],chdata[20],chdata[20:18],
                      chdata[17],chdata[17],chdata[17:15],chdata[14],chdata[14],chdata[14:12],
                      chdata[11],chdata[11],chdata[11:9 ],chdata[8 ],chdata[8 ],chdata[8 :6 ],
                      chdata[5 ],chdata[5 ],chdata[5 :3 ],chdata[2 ],chdata[2 ],chdata[2 :0 ]};
wire [79:0] mtv1_o;
wire [79:0] mtv2_o;
wire [47:0] mtv1_w=(iter_count==5'd0)?47'd0:mtv1;
wire [47:0] mtv2_w=(iter_count==5'd0)?47'd0:mtv2;                                                                                        
wire [79:0]
sumdata1= deca_en ? sumdata1a_o:sumdata1b_o,
sumdata2= deca_en ? sumdata2a_o:sumdata2b_o;
wire [79:0]  sumdata1_w;
wire [79:0]  sumdata2_w;
wire signed [5:0] mtv1_t ={sumdata1[79],sumdata1[79:75]} - {mtv1_w[47],mtv1_w[47],mtv1_w[47],mtv1_w[47:45]};
wire signed [5:0] mtv2_t ={sumdata1[74],sumdata1[74:70]} - {mtv1_w[44],mtv1_w[44],mtv1_w[44],mtv1_w[44:42]};
wire signed [5:0] mtv3_t ={sumdata1[69],sumdata1[69:65]} - {mtv1_w[41],mtv1_w[41],mtv1_w[41],mtv1_w[41:39]};
wire signed [5:0] mtv4_t ={sumdata1[64],sumdata1[64:60]} - {mtv1_w[38],mtv1_w[38],mtv1_w[38],mtv1_w[38:36]};
wire signed [5:0] mtv5_t ={sumdata1[59],sumdata1[59:55]} - {mtv1_w[35],mtv1_w[35],mtv1_w[35],mtv1_w[35:33]};
wire signed [5:0] mtv6_t ={sumdata1[54],sumdata1[54:50]} - {mtv1_w[32],mtv1_w[32],mtv1_w[32],mtv1_w[32:30]};
wire signed [5:0] mtv7_t ={sumdata1[49],sumdata1[49:45]} - {mtv1_w[29],mtv1_w[29],mtv1_w[29],mtv1_w[29:27]};
wire signed [5:0] mtv8_t ={sumdata1[44],sumdata1[44:40]} - {mtv1_w[26],mtv1_w[26],mtv1_w[26],mtv1_w[26:24]};
wire signed [5:0] mtv9_t ={sumdata1[39],sumdata1[39:35]} - {mtv1_w[23],mtv1_w[23],mtv1_w[23],mtv1_w[23:21]};
wire signed [5:0] mtv10_t={sumdata1[34],sumdata1[34:30]} - {mtv1_w[20],mtv1_w[20],mtv1_w[20],mtv1_w[20:18]};
wire signed [5:0] mtv11_t={sumdata1[29],sumdata1[29:25]} - {mtv1_w[17],mtv1_w[17],mtv1_w[17],mtv1_w[17:15]};
wire signed [5:0] mtv12_t={sumdata1[24],sumdata1[24:20]} - {mtv1_w[14],mtv1_w[14],mtv1_w[14],mtv1_w[14:12]};
wire signed [5:0] mtv13_t={sumdata1[19],sumdata1[19:15]} - {mtv1_w[11],mtv1_w[11],mtv1_w[11],mtv1_w[11:9 ]};
wire signed [5:0] mtv14_t={sumdata1[14],sumdata1[14:10]} - {mtv1_w[8 ],mtv1_w[8 ],mtv1_w[8 ],mtv1_w[8 :6 ]};
wire signed [5:0] mtv15_t={sumdata1[9 ],sumdata1[9 :5 ]} - {mtv1_w[5 ],mtv1_w[5 ],mtv1_w[5 ],mtv1_w[5 :3 ]};
wire signed [5:0] mtv16_t={sumdata1[4 ],sumdata1[4 :0 ]} - {mtv1_w[2 ],mtv1_w[2 ],mtv1_w[2 ],mtv1_w[2 :0 ]};

assign mtv1_o[79:75]= (mtv1_t [5] ^ mtv1_t [4]) ? mtv1_t [5] ? {mtv1_t [5],4'b0001} : {mtv1_t [5],4'b1111} : {mtv1_t [5],mtv1_t [3:0]};
assign mtv1_o[74:70]= (mtv2_t [5] ^ mtv2_t [4]) ? mtv2_t [5] ? {mtv2_t [5],4'b0001} : {mtv2_t [5],4'b1111} : {mtv2_t [5],mtv2_t [3:0]};
assign mtv1_o[69:65]= (mtv3_t [5] ^ mtv3_t [4]) ? mtv3_t [5] ? {mtv3_t [5],4'b0001} : {mtv3_t [5],4'b1111} : {mtv3_t [5],mtv3_t [3:0]};
assign mtv1_o[64:60]= (mtv4_t [5] ^ mtv4_t [4]) ? mtv4_t [5] ? {mtv4_t [5],4'b0001} : {mtv4_t [5],4'b1111} : {mtv4_t [5],mtv4_t [3:0]};
assign mtv1_o[59:55]= (mtv5_t [5] ^ mtv5_t [4]) ? mtv5_t [5] ? {mtv5_t [5],4'b0001} : {mtv5_t [5],4'b1111} : {mtv5_t [5],mtv5_t [3:0]};
assign mtv1_o[54:50]= (mtv6_t [5] ^ mtv6_t [4]) ? mtv6_t [5] ? {mtv6_t [5],4'b0001} : {mtv6_t [5],4'b1111} : {mtv6_t [5],mtv6_t [3:0]};
assign mtv1_o[49:45]= (mtv7_t [5] ^ mtv7_t [4]) ? mtv7_t [5] ? {mtv7_t [5],4'b0001} : {mtv7_t [5],4'b1111} : {mtv7_t [5],mtv7_t [3:0]};
assign mtv1_o[44:40]= (mtv8_t [5] ^ mtv8_t [4]) ? mtv8_t [5] ? {mtv8_t [5],4'b0001} : {mtv8_t [5],4'b1111} : {mtv8_t [5],mtv8_t [3:0]};
assign mtv1_o[39:35]= (mtv9_t [5] ^ mtv9_t [4]) ? mtv9_t [5] ? {mtv9_t [5],4'b0001} : {mtv9_t [5],4'b1111} : {mtv9_t [5],mtv9_t [3:0]};
assign mtv1_o[34:30]= (mtv10_t[5] ^ mtv10_t[4]) ? mtv10_t[5] ? {mtv10_t[5],4'b0001} : {mtv10_t[5],4'b1111} : {mtv10_t[5],mtv10_t[3:0]};
assign mtv1_o[29:25]= (mtv11_t[5] ^ mtv11_t[4]) ? mtv11_t[5] ? {mtv11_t[5],4'b0001} : {mtv11_t[5],4'b1111} : {mtv11_t[5],mtv11_t[3:0]};
assign mtv1_o[24:20]= (mtv12_t[5] ^ mtv12_t[4]) ? mtv12_t[5] ? {mtv12_t[5],4'b0001} : {mtv12_t[5],4'b1111} : {mtv12_t[5],mtv12_t[3:0]};
assign mtv1_o[19:15]= (mtv13_t[5] ^ mtv13_t[4]) ? mtv13_t[5] ? {mtv13_t[5],4'b0001} : {mtv13_t[5],4'b1111} : {mtv13_t[5],mtv13_t[3:0]};
assign mtv1_o[14:10]= (mtv14_t[5] ^ mtv14_t[4]) ? mtv14_t[5] ? {mtv14_t[5],4'b0001} : {mtv14_t[5],4'b1111} : {mtv14_t[5],mtv14_t[3:0]};
assign mtv1_o[9 :5 ]= (mtv15_t[5] ^ mtv15_t[4]) ? mtv15_t[5] ? {mtv15_t[5],4'b0001} : {mtv15_t[5],4'b1111} : {mtv15_t[5],mtv15_t[3:0]};
assign mtv1_o[4 :0 ]= (mtv16_t[5] ^ mtv16_t[4]) ? mtv16_t[5] ? {mtv16_t[5],4'b0001} : {mtv16_t[5],4'b1111} : {mtv16_t[5],mtv16_t[3:0]};

wire signed [5:0] mtv17_t={sumdata2[79],sumdata2[79:75]} - {mtv2_w[47],mtv2_w[47],mtv2_w[47],mtv2_w[47:45]};
wire signed [5:0] mtv18_t={sumdata2[74],sumdata2[74:70]} - {mtv2_w[44],mtv2_w[44],mtv2_w[44],mtv2_w[44:42]};
wire signed [5:0] mtv19_t={sumdata2[69],sumdata2[69:65]} - {mtv2_w[41],mtv2_w[41],mtv2_w[41],mtv2_w[41:39]};
wire signed [5:0] mtv20_t={sumdata2[64],sumdata2[64:60]} - {mtv2_w[38],mtv2_w[38],mtv2_w[38],mtv2_w[38:36]};
wire signed [5:0] mtv21_t={sumdata2[59],sumdata2[59:55]} - {mtv2_w[35],mtv2_w[35],mtv2_w[35],mtv2_w[35:33]};
wire signed [5:0] mtv22_t={sumdata2[54],sumdata2[54:50]} - {mtv2_w[32],mtv2_w[32],mtv2_w[32],mtv2_w[32:30]};
wire signed [5:0] mtv23_t={sumdata2[49],sumdata2[49:45]} - {mtv2_w[29],mtv2_w[29],mtv2_w[29],mtv2_w[29:27]};
wire signed [5:0] mtv24_t={sumdata2[44],sumdata2[44:40]} - {mtv2_w[26],mtv2_w[26],mtv2_w[26],mtv2_w[26:24]};
wire signed [5:0] mtv25_t={sumdata2[39],sumdata2[39:35]} - {mtv2_w[23],mtv2_w[23],mtv2_w[23],mtv2_w[23:21]};
wire signed [5:0] mtv26_t={sumdata2[34],sumdata2[34:30]} - {mtv2_w[20],mtv2_w[20],mtv2_w[20],mtv2_w[20:18]};
wire signed [5:0] mtv27_t={sumdata2[29],sumdata2[29:25]} - {mtv2_w[17],mtv2_w[17],mtv2_w[17],mtv2_w[17:15]};
wire signed [5:0] mtv28_t={sumdata2[24],sumdata2[24:20]} - {mtv2_w[14],mtv2_w[14],mtv2_w[14],mtv2_w[14:12]};
wire signed [5:0] mtv29_t={sumdata2[19],sumdata2[19:15]} - {mtv2_w[11],mtv2_w[11],mtv2_w[11],mtv2_w[11:9 ]};
wire signed [5:0] mtv30_t={sumdata2[14],sumdata2[14:10]} - {mtv2_w[8 ],mtv2_w[8 ],mtv2_w[8 ],mtv2_w[8 :6 ]};
wire signed [5:0] mtv31_t={sumdata2[9 ],sumdata2[9 :5 ]} - {mtv2_w[5 ],mtv2_w[5 ],mtv2_w[5 ],mtv2_w[5 :3 ]};
wire signed [5:0] mtv32_t={sumdata2[4 ],sumdata2[4 :0 ]} - {mtv2_w[2 ],mtv2_w[2 ],mtv2_w[2 ],mtv2_w[2 :0 ]};

assign mtv2_o[79:75]= (mtv17_t[5] ^ mtv17_t[4]) ? mtv17_t[5] ? {mtv17_t[5],4'b0001} : {mtv17_t[5],4'b1111} : {mtv17_t[5],mtv17_t[3:0]};
assign mtv2_o[74:70]= (mtv18_t[5] ^ mtv18_t[4]) ? mtv18_t[5] ? {mtv18_t[5],4'b0001} : {mtv18_t[5],4'b1111} : {mtv18_t[5],mtv18_t[3:0]};
assign mtv2_o[69:65]= (mtv19_t[5] ^ mtv19_t[4]) ? mtv19_t[5] ? {mtv19_t[5],4'b0001} : {mtv19_t[5],4'b1111} : {mtv19_t[5],mtv19_t[3:0]};
assign mtv2_o[64:60]= (mtv20_t[5] ^ mtv20_t[4]) ? mtv20_t[5] ? {mtv20_t[5],4'b0001} : {mtv20_t[5],4'b1111} : {mtv20_t[5],mtv20_t[3:0]};
assign mtv2_o[59:55]= (mtv21_t[5] ^ mtv21_t[4]) ? mtv21_t[5] ? {mtv21_t[5],4'b0001} : {mtv21_t[5],4'b1111} : {mtv21_t[5],mtv21_t[3:0]};
assign mtv2_o[54:50]= (mtv22_t[5] ^ mtv22_t[4]) ? mtv22_t[5] ? {mtv22_t[5],4'b0001} : {mtv22_t[5],4'b1111} : {mtv22_t[5],mtv22_t[3:0]};
assign mtv2_o[49:45]= (mtv23_t[5] ^ mtv23_t[4]) ? mtv23_t[5] ? {mtv23_t[5],4'b0001} : {mtv23_t[5],4'b1111} : {mtv23_t[5],mtv23_t[3:0]};
assign mtv2_o[44:40]= (mtv24_t[5] ^ mtv24_t[4]) ? mtv24_t[5] ? {mtv24_t[5],4'b0001} : {mtv24_t[5],4'b1111} : {mtv24_t[5],mtv24_t[3:0]};
assign mtv2_o[39:35]= (mtv25_t[5] ^ mtv25_t[4]) ? mtv25_t[5] ? {mtv25_t[5],4'b0001} : {mtv25_t[5],4'b1111} : {mtv25_t[5],mtv25_t[3:0]};
assign mtv2_o[34:30]= (mtv26_t[5] ^ mtv26_t[4]) ? mtv26_t[5] ? {mtv26_t[5],4'b0001} : {mtv26_t[5],4'b1111} : {mtv26_t[5],mtv26_t[3:0]};
assign mtv2_o[29:25]= (mtv27_t[5] ^ mtv27_t[4]) ? mtv27_t[5] ? {mtv27_t[5],4'b0001} : {mtv27_t[5],4'b1111} : {mtv27_t[5],mtv27_t[3:0]};
assign mtv2_o[24:20]= (mtv28_t[5] ^ mtv28_t[4]) ? mtv28_t[5] ? {mtv28_t[5],4'b0001} : {mtv28_t[5],4'b1111} : {mtv28_t[5],mtv28_t[3:0]};
assign mtv2_o[19:15]= (mtv29_t[5] ^ mtv29_t[4]) ? mtv29_t[5] ? {mtv29_t[5],4'b0001} : {mtv29_t[5],4'b1111} : {mtv29_t[5],mtv29_t[3:0]};
assign mtv2_o[14:10]= (mtv30_t[5] ^ mtv30_t[4]) ? mtv30_t[5] ? {mtv30_t[5],4'b0001} : {mtv30_t[5],4'b1111} : {mtv30_t[5],mtv30_t[3:0]};
assign mtv2_o[9 :5 ]= (mtv31_t[5] ^ mtv31_t[4]) ? mtv31_t[5] ? {mtv31_t[5],4'b0001} : {mtv31_t[5],4'b1111} : {mtv31_t[5],mtv31_t[3:0]};
assign mtv2_o[4 :0 ]= (mtv32_t[5] ^ mtv32_t[4]) ? mtv32_t[5] ? {mtv32_t[5],4'b0001} : {mtv32_t[5],4'b1111} : {mtv32_t[5],mtv32_t[3:0]};


wire signed [5:0] sumdata1_t ={mtv1_o[79],mtv1_o[79:75]} + {ctm1_i[47],ctm1_i[47],ctm1_i[47],ctm1_i[47:45]};
wire signed [5:0] sumdata2_t ={mtv1_o[74],mtv1_o[74:70]} + {ctm1_i[44],ctm1_i[44],ctm1_i[44],ctm1_i[44:42]};
wire signed [5:0] sumdata3_t ={mtv1_o[69],mtv1_o[69:65]} + {ctm1_i[41],ctm1_i[41],ctm1_i[41],ctm1_i[41:39]};
wire signed [5:0] sumdata4_t ={mtv1_o[64],mtv1_o[64:60]} + {ctm1_i[38],ctm1_i[38],ctm1_i[38],ctm1_i[38:36]};
wire signed [5:0] sumdata5_t ={mtv1_o[59],mtv1_o[59:55]} + {ctm1_i[35],ctm1_i[35],ctm1_i[35],ctm1_i[35:33]};
wire signed [5:0] sumdata6_t ={mtv1_o[54],mtv1_o[54:50]} + {ctm1_i[32],ctm1_i[32],ctm1_i[32],ctm1_i[32:30]};
wire signed [5:0] sumdata7_t ={mtv1_o[49],mtv1_o[49:45]} + {ctm1_i[29],ctm1_i[29],ctm1_i[29],ctm1_i[29:27]};
wire signed [5:0] sumdata8_t ={mtv1_o[44],mtv1_o[44:40]} + {ctm1_i[26],ctm1_i[26],ctm1_i[26],ctm1_i[26:24]};
wire signed [5:0] sumdata9_t ={mtv1_o[39],mtv1_o[39:35]} + {ctm1_i[23],ctm1_i[23],ctm1_i[23],ctm1_i[23:21]};
wire signed [5:0] sumdata10_t={mtv1_o[34],mtv1_o[34:30]} + {ctm1_i[20],ctm1_i[20],ctm1_i[20],ctm1_i[20:18]};
wire signed [5:0] sumdata11_t={mtv1_o[29],mtv1_o[29:25]} + {ctm1_i[17],ctm1_i[17],ctm1_i[17],ctm1_i[17:15]};
wire signed [5:0] sumdata12_t={mtv1_o[24],mtv1_o[24:20]} + {ctm1_i[14],ctm1_i[14],ctm1_i[14],ctm1_i[14:12]};
wire signed [5:0] sumdata13_t={mtv1_o[19],mtv1_o[19:15]} + {ctm1_i[11],ctm1_i[11],ctm1_i[11],ctm1_i[11:9 ]};
wire signed [5:0] sumdata14_t={mtv1_o[14],mtv1_o[14:10]} + {ctm1_i[8 ],ctm1_i[8 ],ctm1_i[8 ],ctm1_i[8 :6 ]};
wire signed [5:0] sumdata15_t={mtv1_o[9 ],mtv1_o[9 :5 ]} + {ctm1_i[5 ],ctm1_i[5 ],ctm1_i[5 ],ctm1_i[5 :3 ]};
wire signed [5:0] sumdata16_t={mtv1_o[4 ],mtv1_o[4 :0 ]} + {ctm1_i[2 ],ctm1_i[2 ],ctm1_i[2 ],ctm1_i[2 :0 ]};

assign sumdata1_w[79:75]=(sumdata1_t [5] ^ sumdata1_t [4]) ? sumdata1_t [5] ? {sumdata1_t [5],4'b0001} : {sumdata1_t [5],4'b1111} : {sumdata1_t [5],sumdata1_t [3:0]};
assign sumdata1_w[74:70]=(sumdata2_t [5] ^ sumdata2_t [4]) ? sumdata2_t [5] ? {sumdata2_t [5],4'b0001} : {sumdata2_t [5],4'b1111} : {sumdata2_t [5],sumdata2_t [3:0]};
assign sumdata1_w[69:65]=(sumdata3_t [5] ^ sumdata3_t [4]) ? sumdata3_t [5] ? {sumdata3_t [5],4'b0001} : {sumdata3_t [5],4'b1111} : {sumdata3_t [5],sumdata3_t [3:0]};
assign sumdata1_w[64:60]=(sumdata4_t [5] ^ sumdata4_t [4]) ? sumdata4_t [5] ? {sumdata4_t [5],4'b0001} : {sumdata4_t [5],4'b1111} : {sumdata4_t [5],sumdata4_t [3:0]};
assign sumdata1_w[59:55]=(sumdata5_t [5] ^ sumdata5_t [4]) ? sumdata5_t [5] ? {sumdata5_t [5],4'b0001} : {sumdata5_t [5],4'b1111} : {sumdata5_t [5],sumdata5_t [3:0]};
assign sumdata1_w[54:50]=(sumdata6_t [5] ^ sumdata6_t [4]) ? sumdata6_t [5] ? {sumdata6_t [5],4'b0001} : {sumdata6_t [5],4'b1111} : {sumdata6_t [5],sumdata6_t [3:0]};
assign sumdata1_w[49:45]=(sumdata7_t [5] ^ sumdata7_t [4]) ? sumdata7_t [5] ? {sumdata7_t [5],4'b0001} : {sumdata7_t [5],4'b1111} : {sumdata7_t [5],sumdata7_t [3:0]};
assign sumdata1_w[44:40]=(sumdata8_t [5] ^ sumdata8_t [4]) ? sumdata8_t [5] ? {sumdata8_t [5],4'b0001} : {sumdata8_t [5],4'b1111} : {sumdata8_t [5],sumdata8_t [3:0]};
assign sumdata1_w[39:35]=(sumdata9_t [5] ^ sumdata9_t [4]) ? sumdata9_t [5] ? {sumdata9_t [5],4'b0001} : {sumdata9_t [5],4'b1111} : {sumdata9_t [5],sumdata9_t [3:0]};
assign sumdata1_w[34:30]=(sumdata10_t[5] ^ sumdata10_t[4]) ? sumdata10_t[5] ? {sumdata10_t[5],4'b0001} : {sumdata10_t[5],4'b1111} : {sumdata10_t[5],sumdata10_t[3:0]};
assign sumdata1_w[29:25]=(sumdata11_t[5] ^ sumdata11_t[4]) ? sumdata11_t[5] ? {sumdata11_t[5],4'b0001} : {sumdata11_t[5],4'b1111} : {sumdata11_t[5],sumdata11_t[3:0]};
assign sumdata1_w[24:20]=(sumdata12_t[5] ^ sumdata12_t[4]) ? sumdata12_t[5] ? {sumdata12_t[5],4'b0001} : {sumdata12_t[5],4'b1111} : {sumdata12_t[5],sumdata12_t[3:0]};
assign sumdata1_w[19:15]=(sumdata13_t[5] ^ sumdata13_t[4]) ? sumdata13_t[5] ? {sumdata13_t[5],4'b0001} : {sumdata13_t[5],4'b1111} : {sumdata13_t[5],sumdata13_t[3:0]};
assign sumdata1_w[14:10]=(sumdata14_t[5] ^ sumdata14_t[4]) ? sumdata14_t[5] ? {sumdata14_t[5],4'b0001} : {sumdata14_t[5],4'b1111} : {sumdata14_t[5],sumdata14_t[3:0]};
assign sumdata1_w[9 :5 ]=(sumdata15_t[5] ^ sumdata15_t[4]) ? sumdata15_t[5] ? {sumdata15_t[5],4'b0001} : {sumdata15_t[5],4'b1111} : {sumdata15_t[5],sumdata15_t[3:0]};
assign sumdata1_w[4 :0 ]=(sumdata16_t[5] ^ sumdata16_t[4]) ? sumdata16_t[5] ? {sumdata16_t[5],4'b0001} : {sumdata16_t[5],4'b1111} : {sumdata16_t[5],sumdata16_t[3:0]};

wire signed [5:0] sumdata17_t={mtv2_o[79],mtv2_o[79:75]} + {ctm2_i[47],ctm2_i[47],ctm2_i[47],ctm2_i[47:45]};
wire signed [5:0] sumdata18_t={mtv2_o[74],mtv2_o[74:70]} + {ctm2_i[44],ctm2_i[44],ctm2_i[44],ctm2_i[44:42]};
wire signed [5:0] sumdata19_t={mtv2_o[69],mtv2_o[69:65]} + {ctm2_i[41],ctm2_i[41],ctm2_i[41],ctm2_i[41:39]};
wire signed [5:0] sumdata20_t={mtv2_o[64],mtv2_o[64:60]} + {ctm2_i[38],ctm2_i[38],ctm2_i[38],ctm2_i[38:36]};
wire signed [5:0] sumdata21_t={mtv2_o[59],mtv2_o[59:55]} + {ctm2_i[35],ctm2_i[35],ctm2_i[35],ctm2_i[35:33]};
wire signed [5:0] sumdata22_t={mtv2_o[54],mtv2_o[54:50]} + {ctm2_i[32],ctm2_i[32],ctm2_i[32],ctm2_i[32:30]};
wire signed [5:0] sumdata23_t={mtv2_o[49],mtv2_o[49:45]} + {ctm2_i[29],ctm2_i[29],ctm2_i[29],ctm2_i[29:27]};
wire signed [5:0] sumdata24_t={mtv2_o[44],mtv2_o[44:40]} + {ctm2_i[26],ctm2_i[26],ctm2_i[26],ctm2_i[26:24]};
wire signed [5:0] sumdata25_t={mtv2_o[39],mtv2_o[39:35]} + {ctm2_i[23],ctm2_i[23],ctm2_i[23],ctm2_i[23:21]};
wire signed [5:0] sumdata26_t={mtv2_o[34],mtv2_o[34:30]} + {ctm2_i[20],ctm2_i[20],ctm2_i[20],ctm2_i[20:18]};
wire signed [5:0] sumdata27_t={mtv2_o[29],mtv2_o[29:25]} + {ctm2_i[17],ctm2_i[17],ctm2_i[17],ctm2_i[17:15]};
wire signed [5:0] sumdata28_t={mtv2_o[24],mtv2_o[24:20]} + {ctm2_i[14],ctm2_i[14],ctm2_i[14],ctm2_i[14:12]};
wire signed [5:0] sumdata29_t={mtv2_o[19],mtv2_o[19:15]} + {ctm2_i[11],ctm2_i[11],ctm2_i[11],ctm2_i[11:9 ]};
wire signed [5:0] sumdata30_t={mtv2_o[14],mtv2_o[14:10]} + {ctm2_i[8 ],ctm2_i[8 ],ctm2_i[8 ],ctm2_i[8 :6 ]};
wire signed [5:0] sumdata31_t={mtv2_o[9 ],mtv2_o[9 :5 ]} + {ctm2_i[5 ],ctm2_i[5 ],ctm2_i[5 ],ctm2_i[5 :3 ]};
wire signed [5:0] sumdata32_t={mtv2_o[4 ],mtv2_o[4 :0 ]} + {ctm2_i[2 ],ctm2_i[2 ],ctm2_i[2 ],ctm2_i[2 :0 ]};

assign sumdata2_w[79:75]=(sumdata17_t[5] ^ sumdata17_t[4]) ? sumdata17_t[5] ? {sumdata17_t[5],4'b0001} : {sumdata17_t[5],4'b1111} : {sumdata17_t[5],sumdata17_t[3:0]};
assign sumdata2_w[74:70]=(sumdata18_t[5] ^ sumdata18_t[4]) ? sumdata18_t[5] ? {sumdata18_t[5],4'b0001} : {sumdata18_t[5],4'b1111} : {sumdata18_t[5],sumdata18_t[3:0]};
assign sumdata2_w[69:65]=(sumdata19_t[5] ^ sumdata19_t[4]) ? sumdata19_t[5] ? {sumdata19_t[5],4'b0001} : {sumdata19_t[5],4'b1111} : {sumdata19_t[5],sumdata19_t[3:0]};
assign sumdata2_w[64:60]=(sumdata20_t[5] ^ sumdata20_t[4]) ? sumdata20_t[5] ? {sumdata20_t[5],4'b0001} : {sumdata20_t[5],4'b1111} : {sumdata20_t[5],sumdata20_t[3:0]};
assign sumdata2_w[59:55]=(sumdata21_t[5] ^ sumdata21_t[4]) ? sumdata21_t[5] ? {sumdata21_t[5],4'b0001} : {sumdata21_t[5],4'b1111} : {sumdata21_t[5],sumdata21_t[3:0]};
assign sumdata2_w[54:50]=(sumdata22_t[5] ^ sumdata22_t[4]) ? sumdata22_t[5] ? {sumdata22_t[5],4'b0001} : {sumdata22_t[5],4'b1111} : {sumdata22_t[5],sumdata22_t[3:0]};
assign sumdata2_w[49:45]=(sumdata23_t[5] ^ sumdata23_t[4]) ? sumdata23_t[5] ? {sumdata23_t[5],4'b0001} : {sumdata23_t[5],4'b1111} : {sumdata23_t[5],sumdata23_t[3:0]};
assign sumdata2_w[44:40]=(sumdata24_t[5] ^ sumdata24_t[4]) ? sumdata24_t[5] ? {sumdata24_t[5],4'b0001} : {sumdata24_t[5],4'b1111} : {sumdata24_t[5],sumdata24_t[3:0]};
assign sumdata2_w[39:35]=(sumdata25_t[5] ^ sumdata25_t[4]) ? sumdata25_t[5] ? {sumdata25_t[5],4'b0001} : {sumdata25_t[5],4'b1111} : {sumdata25_t[5],sumdata25_t[3:0]};
assign sumdata2_w[34:30]=(sumdata26_t[5] ^ sumdata26_t[4]) ? sumdata26_t[5] ? {sumdata26_t[5],4'b0001} : {sumdata26_t[5],4'b1111} : {sumdata26_t[5],sumdata26_t[3:0]};
assign sumdata2_w[29:25]=(sumdata27_t[5] ^ sumdata27_t[4]) ? sumdata27_t[5] ? {sumdata27_t[5],4'b0001} : {sumdata27_t[5],4'b1111} : {sumdata27_t[5],sumdata27_t[3:0]};
assign sumdata2_w[24:20]=(sumdata28_t[5] ^ sumdata28_t[4]) ? sumdata28_t[5] ? {sumdata28_t[5],4'b0001} : {sumdata28_t[5],4'b1111} : {sumdata28_t[5],sumdata28_t[3:0]};
assign sumdata2_w[19:15]=(sumdata29_t[5] ^ sumdata29_t[4]) ? sumdata29_t[5] ? {sumdata29_t[5],4'b0001} : {sumdata29_t[5],4'b1111} : {sumdata29_t[5],sumdata29_t[3:0]};
assign sumdata2_w[14:10]=(sumdata30_t[5] ^ sumdata30_t[4]) ? sumdata30_t[5] ? {sumdata30_t[5],4'b0001} : {sumdata30_t[5],4'b1111} : {sumdata30_t[5],sumdata30_t[3:0]};
assign sumdata2_w[9 :5 ]=(sumdata31_t[5] ^ sumdata31_t[4]) ? sumdata31_t[5] ? {sumdata31_t[5],4'b0001} : {sumdata31_t[5],4'b1111} : {sumdata31_t[5],sumdata31_t[3:0]};
assign sumdata2_w[4 :0 ]=(sumdata32_t[5] ^ sumdata32_t[4]) ? sumdata32_t[5] ? {sumdata32_t[5],4'b0001} : {sumdata32_t[5],4'b1111} : {sumdata32_t[5],sumdata32_t[3:0]};

wire [79:0]
   sumdata1_a=(data_wrsa)?chdata_w:sumdata1_w,
   sumdata2_a=(data_wrsa)?chdata_w:sumdata2_w,
   sumdata1_b=(data_wrsb)?chdata_w:sumdata1_w,
   sumdata2_b=(data_wrsb)?chdata_w:sumdata2_w;

memblock64x80 mem1_a(
           .A(addrcha1_w),
         .CEN(mema_en),
         .CLK(CLK),
         .D(sumdata1_a),
         .WEN(chmemwra1_en),
         .Q(sumdata1a_o)
         );
memblock64x80 mem2_a(
           .A(addrcha2_w),
         .CEN(mema_en),
         .CLK(CLK),
         .D(sumdata2_a),
         .WEN(chmemwra2_en),
         .Q(sumdata2a_o)
         );
memblock64x80 mem1_b(
           .A(addrchb1_w),
         .CEN(memb_en),
         .CLK(CLK),
         .D(sumdata1_b),
         .WEN(chmemwrb1_en),
         .Q(sumdata1b_o)
         );
memblock64x80 mem2_b(
           .A(addrchb2_w),
         .CEN(memb_en),
         .CLK(CLK),
         .D(sumdata2_b),
         .WEN(chmemwrb2_en),
         .Q(sumdata2b_o)
         );

assign addr1a_w= (section==2'b00)? {layer_i,section,addr_count1_1}:
                 (section==2'b01)? {layer_i,section,addr_count1_2}:
                 (section==2'b10)? {layer_i,section,addr_count1_3}:
                                   {layer_i,section,addr_count1_4};
assign addr2a_w= (section==2'b00)? {layer_i,section,addr_count2_1}:
                 (section==2'b01)? {layer_i,section,addr_count2_2}:
                 (section==2'b10)? {layer_i,section,addr_count2_3}:
                                   {layer_i,section,addr_count2_4};

wire [16:1] sgn;
wire keep_min=(vncn_count>4'd4);

wire [95:0] vtc;
wire [2:0] vtc1_1 =vtc[ 2: 0];
wire [2:0] vtc2_1 =vtc[ 5: 3];
wire [2:0] vtc1_2 =vtc[ 8: 6];
wire [2:0] vtc2_2 =vtc[11: 9];
wire [2:0] vtc1_3 =vtc[14:12];
wire [2:0] vtc2_3 =vtc[17:15];
wire [2:0] vtc1_4 =vtc[20:18];
wire [2:0] vtc2_4 =vtc[23:21];
wire [2:0] vtc1_5 =vtc[26:24];
wire [2:0] vtc2_5 =vtc[29:27];
wire [2:0] vtc1_6 =vtc[32:30];
wire [2:0] vtc2_6 =vtc[35:33];
wire [2:0] vtc1_7 =vtc[38:36];
wire [2:0] vtc2_7 =vtc[41:39];
wire [2:0] vtc1_8 =vtc[44:42];
wire [2:0] vtc2_8 =vtc[47:45];
wire [2:0] vtc1_9 =vtc[50:48];
wire [2:0] vtc2_9 =vtc[53:51];
wire [2:0] vtc1_10=vtc[56:54];
wire [2:0] vtc2_10=vtc[59:57];
wire [2:0] vtc1_11=vtc[62:60];
wire [2:0] vtc2_11=vtc[65:63];
wire [2:0] vtc1_12=vtc[68:66];
wire [2:0] vtc2_12=vtc[71:69];
wire [2:0] vtc1_13=vtc[74:72];
wire [2:0] vtc2_13=vtc[77:75];
wire [2:0] vtc1_14=vtc[80:78];
wire [2:0] vtc2_14=vtc[83:81];
wire [2:0] vtc1_15=vtc[86:84];
wire [2:0] vtc2_15=vtc[89:87];
wire [2:0] vtc1_16=vtc[92:90];
wire [2:0] vtc2_16=vtc[95:93];

CNP CNP1(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[1]),.keep_min(keep_min),
         .min_r(min_i1),.secmin_r(secmin_i1),
         .min_loc(min_loc[1]),
         .vtc_1(vtc1_1),.vtc_2(vtc2_1),
         .ctm_1(ctm1_1),.ctm_2(ctm2_1),
         .min(min1),.sgn(sgn[1])
        );
CNP CNP2(
         .CLK(CLK), .RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[2]),.keep_min(keep_min),
         .min_r(min_i2),.secmin_r(secmin_i2),
         .min_loc(min_loc[2]),
         .vtc_1(vtc1_2),.vtc_2(vtc2_2),
         .ctm_1(ctm1_2),.ctm_2(ctm2_2),
         .min(min2),.sgn(sgn[2])
        );
CNP CNP3(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[3]),.keep_min(keep_min),
         .min_r(min_i3),.secmin_r(secmin_i3),
         .min_loc(min_loc[3]),
         .vtc_1(vtc1_3),.vtc_2(vtc2_3),
         .ctm_1(ctm1_3),.ctm_2(ctm2_3),
         .min(min3),.sgn(sgn[3])
        );
CNP CNP4(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[4]),.keep_min(keep_min),
         .min_r(min_i4),.secmin_r(secmin_i4),
         .min_loc(min_loc[4]),
         .vtc_1(vtc1_4),.vtc_2(vtc2_4),
         .ctm_1(ctm1_4),.ctm_2(ctm2_4),
         .min(min4),.sgn(sgn[4])
        );
CNP CNP5(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[5]),.keep_min(keep_min),
         .min_r(min_i5),.secmin_r(secmin_i5),
         .min_loc(min_loc[5]),
         .vtc_1(vtc1_5),.vtc_2(vtc2_5),
         .ctm_1(ctm1_5),.ctm_2(ctm2_5),
         .min(min5),.sgn(sgn[5])
        );
CNP CNP6(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[6]),.keep_min(keep_min),
         .min_r(min_i6),.secmin_r(secmin_i6),
         .min_loc(min_loc[6]),
         .vtc_1(vtc1_6),.vtc_2(vtc2_6),
         .ctm_1(ctm1_6),.ctm_2(ctm2_6),
         .min(min6),.sgn(sgn[6])
        );
CNP CNP7(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[7]),.keep_min(keep_min),
         .min_r(min_i7),.secmin_r(secmin_i7),
         .min_loc(min_loc[7]),
         .vtc_1(vtc1_7),.vtc_2(vtc2_7),
         .ctm_1(ctm1_7),.ctm_2(ctm2_7),
         .min(min7),.sgn(sgn[7])
        );
CNP CNP8(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[8]),.keep_min(keep_min),
         .min_r(min_i8),.secmin_r(secmin_i8),
         .min_loc(min_loc[8]),
         .vtc_1(vtc1_8),.vtc_2(vtc2_8),
         .ctm_1(ctm1_8),.ctm_2(ctm2_8),
         .min(min8),.sgn(sgn[8])
        );
CNP CNP9(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[9]),.keep_min(keep_min),
         .min_r(min_i9),.secmin_r(secmin_i9),
         .min_loc(min_loc[9]),
         .vtc_1(vtc1_9),.vtc_2(vtc2_9),
         .ctm_1(ctm1_9),.ctm_2(ctm2_9),
         .min(min9),.sgn(sgn[9])
        );
CNP CNP10(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[10]),.keep_min(keep_min),
         .min_r(min_i10),.secmin_r(secmin_i10),
         .min_loc(min_loc[10]),
         .vtc_1(vtc1_10),.vtc_2(vtc2_10),
         .ctm_1(ctm1_10),.ctm_2(ctm2_10),
         .min(min10),.sgn(sgn[10])
        );
CNP CNP11(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[11]),.keep_min(keep_min),
         .min_r(min_i11),.secmin_r(secmin_i11),
         .min_loc(min_loc[11]),
         .vtc_1(vtc1_11),.vtc_2(vtc2_11),
         .ctm_1(ctm1_11),.ctm_2(ctm2_11),
         .min(min11),.sgn(sgn[11])
        );
CNP CNP12(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[12]),.keep_min(keep_min),
         .min_r(min_i12),.secmin_r(secmin_i12),
         .min_loc(min_loc[12]),
         .vtc_1(vtc1_12),.vtc_2(vtc2_12),
         .ctm_1(ctm1_12),.ctm_2(ctm2_12),
         .min(min12),.sgn(sgn[12])
        );
CNP CNP13(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[13]),.keep_min(keep_min),
         .min_r(min_i13),.secmin_r(secmin_i13),
         .min_loc(min_loc[13]),
         .vtc_1(vtc1_13),.vtc_2(vtc2_13),
         .ctm_1(ctm1_13),.ctm_2(ctm2_13),
         .min(min13),.sgn(sgn[13])
        );
CNP CNP14(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[14]),.keep_min(keep_min),
         .min_r(min_i14),.secmin_r(secmin_i14),
         .min_loc(min_loc[14]),
         .vtc_1(vtc1_14),.vtc_2(vtc2_14),
         .ctm_1(ctm1_14),.ctm_2(ctm2_14),
         .min(min14),.sgn(sgn[14])
        );
CNP CNP15(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[15]),.keep_min(keep_min),
         .min_r(min_i15),.secmin_r(secmin_i15),
         .min_loc(min_loc[15]),
         .vtc_1(vtc1_15),.vtc_2(vtc2_15),
         .ctm_1(ctm1_15),.ctm_2(ctm2_15),
         .min(min15),.sgn(sgn[15])
        );
CNP CNP16(
         .CLK(CLK),.RESET_N(RESET_N),
         .vncn_en(vncn_en),.section(section_r),
         .totsgn(sgn_i[16]),.keep_min(keep_min),
         .min_r(min_i16),.secmin_r(secmin_i16),
         .min_loc(min_loc[16]),
         .vtc_1(vtc1_16),.vtc_2(vtc2_16),
         .ctm_1(ctm1_16),.ctm_2(ctm2_16),
         .min(min16),.sgn(sgn[16])
        );

wire [47:0]
  ctm1 ={ctm1_16,ctm1_15,ctm1_14,ctm1_13,
         ctm1_12,ctm1_11,ctm1_10,ctm1_9,
         ctm1_8,ctm1_7,ctm1_6,ctm1_5,
         ctm1_4,ctm1_3,ctm1_2,ctm1_1},
  ctm2 ={ctm2_16,ctm2_15,ctm2_14,ctm2_13,
         ctm2_12,ctm2_11,ctm2_10,ctm2_9,
         ctm2_8,ctm2_7,ctm2_6,ctm2_5,
         ctm2_4,ctm2_3,ctm2_2,ctm2_1};

wire [47:0] rtm1a_w =ctm1_i;
wire [47:0] rtm2a_w =ctm2_i;


wire memwr_en =deca_en ? memwra_en:memwrb_en;
wire mem_en= dec_en ;

memblock256x48 mem1(
         .A(addr1a_w),
         .CEN(mem_en),
         .CLK(CLK),
         .D(rtm1a_w),
         .WEN(memwr_en),
         .Q(mtv1)
         );
memblock256x48 mem2(
         .A(addr2a_w),
         .CEN(mem_en),
         .CLK(CLK),
         .D(rtm2a_w),
         .WEN(memwr_en),
         .Q(mtv2)
         );

VNPgroup VNPgroup(
                  .stv1_w (mtv1_i ), .stv2_w (mtv2_i ),
                  .summtv1_w  (sumdata1_i ), .summtv2_w  (sumdata2_i ),
                  .hardbit(sr_hb),
                  .vtc(vtc));
endmodule

module VNPgroup(
                stv1_w,stv2_w,
                summtv1_w,summtv2_w,
                hardbit,
                vtc);

input  [79:0] stv1_w,stv2_w;
input  [79:0] summtv1_w,summtv2_w;
output [31:0] hardbit;
output [95:0] vtc;

wire signed [4:0] sumout1 =stv1_w[4:0]  ;
wire signed [4:0] sumout2 =stv2_w[4:0]  ;
wire signed [4:0] sumout3 =stv1_w[9:5]  ;
wire signed [4:0] sumout4 =stv2_w[9:5]  ;
wire signed [4:0] sumout5 =stv1_w[14:10] ;
wire signed [4:0] sumout6 =stv2_w[14:10] ;
wire signed [4:0] sumout7 =stv1_w[19:15];
wire signed [4:0] sumout8 =stv2_w[19:15];
wire signed [4:0] sumout9 =stv1_w[24:20];
wire signed [4:0] sumout10=stv2_w[24:20];
wire signed [4:0] sumout11=stv1_w[29:25];
wire signed [4:0] sumout12=stv2_w[29:25];
wire signed [4:0] sumout13=stv1_w[34:30];
wire signed [4:0] sumout14=stv2_w[34:30];
wire signed [4:0] sumout15=stv1_w[39:35];
wire signed [4:0] sumout16=stv2_w[39:35];
wire signed [4:0] sumout17=stv1_w[44:40];
wire signed [4:0] sumout18=stv2_w[44:40];
wire signed [4:0] sumout19=stv1_w[49:45];
wire signed [4:0] sumout20=stv2_w[49:45];
wire signed [4:0] sumout21=stv1_w[54:50];
wire signed [4:0] sumout22=stv2_w[54:50];
wire signed [4:0] sumout23=stv1_w[59:55];
wire signed [4:0] sumout24=stv2_w[59:55];
wire signed [4:0] sumout25=stv1_w[64:60];
wire signed [4:0] sumout26=stv2_w[64:60];
wire signed [4:0] sumout27=stv1_w[69:65];
wire signed [4:0] sumout28=stv2_w[69:65];
wire signed [4:0] sumout29=stv1_w[74:70];
wire signed [4:0] sumout30=stv2_w[74:70];
wire signed [4:0] sumout31=stv1_w[79:75];
wire signed [4:0] sumout32=stv2_w[79:75];
wire signed [4:0] summtv1 =summtv1_w[4:0]  ;
wire signed [4:0] summtv2 =summtv2_w[4:0]  ;
wire signed [4:0] summtv3 =summtv1_w[9:5]  ;
wire signed [4:0] summtv4 =summtv2_w[9:5]  ;
wire signed [4:0] summtv5 =summtv1_w[14:10] ;
wire signed [4:0] summtv6 =summtv2_w[14:10] ;
wire signed [4:0] summtv7 =summtv1_w[19:15];
wire signed [4:0] summtv8 =summtv2_w[19:15];
wire signed [4:0] summtv9 =summtv1_w[24:20];
wire signed [4:0] summtv10=summtv2_w[24:20];
wire signed [4:0] summtv11=summtv1_w[29:25];
wire signed [4:0] summtv12=summtv2_w[29:25];
wire signed [4:0] summtv13=summtv1_w[34:30];
wire signed [4:0] summtv14=summtv2_w[34:30];
wire signed [4:0] summtv15=summtv1_w[39:35];
wire signed [4:0] summtv16=summtv2_w[39:35];
wire signed [4:0] summtv17=summtv1_w[44:40];
wire signed [4:0] summtv18=summtv2_w[44:40];
wire signed [4:0] summtv19=summtv1_w[49:45];
wire signed [4:0] summtv20=summtv2_w[49:45];
wire signed [4:0] summtv21=summtv1_w[54:50];
wire signed [4:0] summtv22=summtv2_w[54:50];
wire signed [4:0] summtv23=summtv1_w[59:55];
wire signed [4:0] summtv24=summtv2_w[59:55];
wire signed [4:0] summtv25=summtv1_w[64:60];
wire signed [4:0] summtv26=summtv2_w[64:60];
wire signed [4:0] summtv27=summtv1_w[69:65];
wire signed [4:0] summtv28=summtv2_w[69:65];
wire signed [4:0] summtv29=summtv1_w[74:70];
wire signed [4:0] summtv30=summtv2_w[74:70];
wire signed [4:0] summtv31=summtv1_w[79:75];
wire signed [4:0] summtv32=summtv2_w[79:75];
//VNP1

wire signed [2:0] vtc1=( (sumout1[3] ^  sumout1[4]) |
                         (sumout1[2] ^  sumout1[4]) ) ?
                         (sumout1[4])?{sumout1[4],2'b01}:{sumout1[4],2'b11}:
                         {sumout1[4],sumout1[1:0]};
//VNP2

wire signed [2:0] vtc2=( (sumout2[3] ^  sumout2[4]) |
                         (sumout2[2] ^  sumout2[4]) ) ?
                        (sumout2[4])?{sumout2[4],2'b01}:{sumout2[4],2'b11}:
                        {sumout2[4],sumout2[1:0]};
//VNP3

wire signed [2:0] vtc3=( (sumout3[3] ^  sumout3[4]) |
                         (sumout3[2] ^  sumout3[4]) ) ?
                        (sumout3[4])?{sumout3[4],2'b01}:{sumout3[4],2'b11}:
                        {sumout3[4],sumout3[1:0]};
//VNP4

wire signed [2:0] vtc4=( (sumout4[3] ^  sumout4[4]) |
                         (sumout4[2] ^  sumout4[4]) ) ?
                        (sumout4[4])?{sumout4[4],2'b01}:{sumout4[4],2'b11}:
                        {sumout4[4],sumout4[1:0]};
//VNP5

wire signed [2:0] vtc5=( (sumout5[3] ^  sumout5[4]) |
                         (sumout5[2] ^  sumout5[4]) ) ?
                        (sumout5[4])?{sumout5[4],2'b01}:{sumout5[4],2'b11}:
                        {sumout5[4],sumout5[1:0]};
//VNP6

wire signed [2:0] vtc6=( (sumout6[3] ^  sumout6[4]) |
                         (sumout6[2] ^  sumout6[4]) ) ?
                        (sumout6[4])?{sumout6[4],2'b01}:{sumout6[4],2'b11}:
                        {sumout6[4],sumout6[1:0]};
//VNP7

wire signed [2:0] vtc7=( (sumout7[3] ^  sumout7[4]) |
                         (sumout7[2] ^  sumout7[4]) ) ?
                        (sumout7[4])?{sumout7[4],2'b01}:{sumout7[4],2'b11}:
                        {sumout7[4],sumout7[1:0]};
//VNP8

wire signed [2:0] vtc8=( (sumout8[3] ^  sumout8[4]) |
                         (sumout8[2] ^  sumout8[4]) ) ?
                        (sumout8[4])?{sumout8[4],2'b01}:{sumout8[4],2'b11}:
                        {sumout8[4],sumout8[1:0]};
//VNP9

wire signed [2:0] vtc9=( (sumout9[3] ^  sumout9[4]) |
                         (sumout9[2] ^  sumout9[4]) ) ?
                        (sumout9[4])?{sumout9[4],2'b01}:{sumout9[4],2'b11}:
                        {sumout9[4],sumout9[1:0]};
//VNP10

wire signed [2:0] vtc10=( (sumout10[3] ^  sumout10[4]) |
                          (sumout10[2] ^  sumout10[4]) ) ?
                         (sumout10[4])?{sumout10[4],2'b01}:{sumout10[4],2'b11}:
                         {sumout10[4],sumout10[1:0]};
//VNP11

wire signed [2:0] vtc11=( (sumout11[3] ^  sumout11[4]) |
                          (sumout11[2] ^  sumout11[4]) ) ?
                         (sumout11[4])?{sumout11[4],2'b01}:{sumout11[4],2'b11}:
                         {sumout11[4],sumout11[1:0]};
//VNP12

wire signed [2:0] vtc12=( (sumout12[3] ^  sumout12[4]) |
                          (sumout12[2] ^  sumout12[4]) ) ?
                         (sumout12[4])?{sumout12[4],2'b01}:{sumout12[4],2'b11}:
                         {sumout12[4],sumout12[1:0]};
//VNP13

wire signed [2:0] vtc13=( (sumout13[3] ^  sumout13[4]) |
                          (sumout13[2] ^  sumout13[4]) ) ?
                         (sumout13[4])?{sumout13[4],2'b01}:{sumout13[4],2'b11}:
                         {sumout13[4],sumout13[1:0]};
//VNP14

wire signed [2:0] vtc14=( (sumout14[3] ^  sumout14[4]) |
                          (sumout14[2] ^  sumout14[4]) ) ?
                         (sumout14[4])?{sumout14[4],2'b01}:{sumout14[4],2'b11}:
                         {sumout14[4],sumout14[1:0]};
//VNP15

wire signed [2:0] vtc15=( (sumout15[3] ^  sumout15[4]) |
                          (sumout15[2] ^  sumout15[4]) ) ?
                         (sumout15[4])?{sumout15[4],2'b01}:{sumout15[4],2'b11}:
                         {sumout15[4],sumout15[1:0]};
//VNP16

wire signed [2:0] vtc16=( (sumout16[3] ^  sumout16[4]) |
                          (sumout16[2] ^  sumout16[4]) ) ?
                         (sumout16[4])?{sumout16[4],2'b01}:{sumout16[4],2'b11}:
                         {sumout16[4],sumout16[1:0]};
//VNP17

wire signed [2:0] vtc17=( (sumout17[3] ^  sumout17[4]) |
                          (sumout17[2] ^  sumout17[4]) ) ?
                         (sumout17[4])?{sumout17[4],2'b01}:{sumout17[4],2'b11}:
                         {sumout17[4],sumout17[1:0]};
//VNP18

wire signed [2:0] vtc18=( (sumout18[3] ^  sumout18[4]) |
                          (sumout18[2] ^  sumout18[4]) ) ?
                         (sumout18[4])?{sumout18[4],2'b01}:{sumout18[4],2'b11}:
                         {sumout18[4],sumout18[1:0]};
//VNP19

wire signed [2:0] vtc19=( (sumout19[3] ^  sumout19[4]) |
                          (sumout19[2] ^  sumout19[4]) ) ?
                         (sumout19[4])?{sumout19[4],2'b01}:{sumout19[4],2'b11}:
                         {sumout19[4],sumout19[1:0]};
//VNP20

wire signed [2:0] vtc20=( (sumout20[3] ^  sumout20[4]) |
                          (sumout20[2] ^  sumout20[4]) ) ?
                         (sumout20[4])?{sumout20[4],2'b01}:{sumout20[4],2'b11}:
                         {sumout20[4],sumout20[1:0]};
//VNP21

wire signed [2:0] vtc21=( (sumout21[3] ^  sumout21[4]) |
                          (sumout21[2] ^  sumout21[4]) ) ?
                         (sumout21[4])?{sumout21[4],2'b01}:{sumout21[4],2'b11}:
                         {sumout21[4],sumout21[1:0]};
//VNP22

wire signed [2:0] vtc22=( (sumout22[3] ^  sumout22[4]) |
                          (sumout22[2] ^  sumout22[4]) ) ?
                         (sumout22[4])?{sumout22[4],2'b01}:{sumout22[4],2'b11}:
                         {sumout22[4],sumout22[1:0]};
//VNP23

wire signed [2:0] vtc23=( (sumout23[3] ^  sumout23[4]) |
                          (sumout23[2] ^  sumout23[4]) ) ?
                         (sumout23[4])?{sumout23[4],2'b01}:{sumout23[4],2'b11}:
                         {sumout23[4],sumout23[1:0]};
//VNP24

wire signed [2:0] vtc24=( (sumout24[3] ^  sumout24[4]) |
                          (sumout24[2] ^  sumout24[4]) ) ?
                         (sumout24[4])?{sumout24[4],2'b01}:{sumout24[4],2'b11}:
                         {sumout24[4],sumout24[1:0]};
//VNP25
wire signed [2:0] vtc25=( (sumout25[3] ^  sumout25[4]) |
                          (sumout25[2] ^  sumout25[4]) ) ?
                         (sumout25[4])?{sumout25[4],2'b01}:{sumout25[4],2'b11}:
                         {sumout25[4],sumout25[1:0]};
//VNP26

wire signed [2:0] vtc26=( (sumout26[3] ^  sumout26[4]) |
                          (sumout26[2] ^  sumout26[4]) ) ?
                         (sumout26[4])?{sumout26[4],2'b01}:{sumout26[4],2'b11}:
                         {sumout26[4],sumout26[1:0]};
//VNP27
wire signed [2:0] vtc27=(((~sumout27[2] | ~sumout27[3]) &  sumout27[4]) |
                         (( sumout27[2] |  sumout27[3]) & ~sumout27[4]))?
                         (sumout27[4])?{sumout27[4],2'b01}:{sumout27[4],2'b11}:
                         {sumout27[4],sumout27[1:0]};
//VNP28

wire signed [2:0] vtc28=( (sumout28[3] ^  sumout28[4]) |
                          (sumout28[2] ^  sumout28[4]) ) ?
                         (sumout28[4])?{sumout28[4],2'b01}:{sumout28[4],2'b11}:
                         {sumout28[4],sumout28[1:0]};
//VNP29
wire signed [2:0] vtc29=( (sumout29[3] ^  sumout29[4]) |
                          (sumout29[2] ^  sumout29[4]) ) ?
                         (sumout29[4])?{sumout29[4],2'b01}:{sumout29[4],2'b11}:
                         {sumout29[4],sumout29[1:0]};
//VNP30

wire signed [2:0] vtc30=( (sumout30[3] ^  sumout30[4]) |
                          (sumout30[2] ^  sumout30[4]) ) ?
                         (sumout30[4])?{sumout30[4],2'b01}:{sumout30[4],2'b11}:
                         {sumout30[4],sumout30[1:0]};
//VNP31

wire signed [2:0] vtc31=( (sumout31[3] ^  sumout31[4]) |
                          (sumout31[2] ^  sumout31[4]) ) ?
                         (sumout31[4])?{sumout31[4],2'b01}:{sumout31[4],2'b11}:
                         {sumout31[4],sumout31[1:0]};
//VNP32

wire signed [2:0] vtc32=( (sumout32[3] ^  sumout32[4]) |
                          (sumout32[2] ^  sumout32[4]) ) ?
                         (sumout32[4])?{sumout32[4],2'b01}:{sumout32[4],2'b11}:
                         {sumout32[4],sumout32[1:0]};


wire [95:0] vtc={vtc32,vtc31,vtc30,vtc29,
                 vtc28,vtc27,vtc26,vtc25,
                 vtc24,vtc23,vtc22,vtc21,
                 vtc20,vtc19,vtc18,vtc17,
                 vtc16,vtc15,vtc14,vtc13,
                 vtc12,vtc11,vtc10,vtc9,
                 vtc8,vtc7,vtc6,vtc5,
                 vtc4,vtc3,vtc2,vtc1};

wire [31:0] hardbit={summtv2 [4], summtv4 [4],  summtv6 [4],  summtv8 [4],
                     summtv10[4], summtv12 [4], summtv14 [4], summtv16[4],
                     summtv18[4], summtv20 [4], summtv22[4],  summtv24[4],
                     summtv26[4], summtv28 [4], summtv30[4],  summtv32[4],
                     summtv1 [4], summtv3 [4],  summtv5[4],   summtv7 [4],
                     summtv9 [4], summtv11[4],  summtv13[4],  summtv15[4],
                     summtv17[4], summtv19 [4], summtv21[4],  summtv23[4],
                     summtv25[4], summtv27 [4], summtv29[4],  summtv31[4]};
endmodule
module  rotatreg(
                 CLK,RESET_N,
                 load_data_en,start_Ldata,
                 data_wrsa,data_wrsb,
                 chdata,
                      chdata_o,
                 memid,memgroup,section_ch);

input CLK,RESET_N, load_data_en,start_Ldata,
      data_wrsa,data_wrsb;
input [47:0] chdata;
output [47:0] chdata_o;
output [2:0] memid;
output [2:0] memgroup;
output [1:0] section_ch;
reg [1:0] section_ch;
reg [4:0] counter;
reg [2:0] memid;
reg [2:0] memgroup;
reg [47:0] chdata_r1 [0:15];
reg [47:0] chdata_r2 [0:15];
reg [47:0] chdata_o;
wire [47:0] chdata_w;

assign
  chdata_w[2 :0] =(chdata[2 ])?
                  {chdata[2 ],~chdata[1:0]+2'd1}:chdata[2:0],
  chdata_w[5 :3] =(chdata[5 ])?
                  {chdata[5 ],~chdata[4:3]+2'd1}:chdata[5:3],
  chdata_w[8 :6] =(chdata[8 ])?
                  {chdata[8 ],~chdata[7:6]+2'd1}:chdata[8:6],
  chdata_w[11:9] =(chdata[11])?
                  {chdata[11],~chdata[10:9]+2'd1}:chdata[11:9],
  chdata_w[14:12]=(chdata[14])?
                  {chdata[14],~chdata[13:12]+2'd1}:chdata[14:12],
  chdata_w[17:15]=(chdata[17])?
                  {chdata[17],~chdata[16:15]+2'd1}:chdata[17:15],
  chdata_w[20:18]=(chdata[20])?
                  {chdata[20],~chdata[19:18]+2'd1}:chdata[20:18],
  chdata_w[23:21]=(chdata[23])?
                  {chdata[23],~chdata[22:21]+2'd1}:chdata[23:21],
  chdata_w[26:24]=(chdata[26])?
                  {chdata[26],~chdata[25:24]+2'd1}:chdata[26:24],
  chdata_w[29:27]=(chdata[29])?
                  {chdata[29],~chdata[28:27]+2'd1}:chdata[29:27],
  chdata_w[32:30]=(chdata[32])?
                  {chdata[32],~chdata[31:30]+2'd1}:chdata[32:30],
  chdata_w[35:33]=(chdata[35])?
                  {chdata[35],~chdata[34:33]+2'd1}:chdata[35:33],
  chdata_w[38:36]=(chdata[38])?
                  {chdata[38],~chdata[37:36]+2'd1}:chdata[38:36],
  chdata_w[41:39]=(chdata[41])?
                  {chdata[41],~chdata[40:39]+2'd1}:chdata[41:39],
  chdata_w[44:42]=(chdata[44])?
                  {chdata[44],~chdata[43:42]+2'd1}:chdata[44:42],
  chdata_w[47:45]=(chdata[47])?
                  {chdata[47],~chdata[46:45]+2'd1}:chdata[47:45];

always @(*)
begin
  case(counter)
    5'd 0:chdata_o={chdata_r2[0 ][ 2: 0],chdata_r2[1 ][ 2: 0],
                     chdata_r2[2 ][ 2: 0],chdata_r2[3 ][ 2: 0],
                     chdata_r2[4 ][ 2: 0],chdata_r2[5 ][ 2: 0],
                     chdata_r2[6 ][ 2: 0],chdata_r2[7 ][ 2: 0],
                     chdata_r2[8 ][ 2: 0],chdata_r2[9 ][ 2: 0],
                     chdata_r2[10 ][ 2: 0],chdata_r2[11 ][ 2: 0],
                     chdata_r2[12 ][ 2: 0],chdata_r2[13 ][ 2: 0],
                     chdata_r2[14 ][ 2: 0],chdata_r2[15][ 2: 0]};
    5'd 1:chdata_o={chdata_r2[0 ][ 5: 3],chdata_r2[1 ][ 5: 3],
                     chdata_r2[2 ][ 5: 3],chdata_r2[3 ][ 5: 3],
                     chdata_r2[4 ][ 5: 3],chdata_r2[5 ][ 5: 3],
                     chdata_r2[6 ][ 5: 3],chdata_r2[7 ][ 5: 3],
                     chdata_r2[8 ][ 5: 3],chdata_r2[9 ][ 5: 3],
                     chdata_r2[10 ][ 5: 3],chdata_r2[11 ][ 5: 3],
                     chdata_r2[12 ][ 5: 3],chdata_r2[13 ][ 5: 3],
                     chdata_r2[14 ][ 5: 3],chdata_r2[15][ 5: 3]};
    5'd 2:chdata_o={chdata_r2[0 ][ 8: 6],chdata_r2[1 ][ 8: 6],
                     chdata_r2[2 ][ 8: 6],chdata_r2[3 ][ 8: 6],
                     chdata_r2[4 ][ 8: 6],chdata_r2[5 ][ 8: 6],
                     chdata_r2[6 ][ 8: 6],chdata_r2[7 ][ 8: 6],
                     chdata_r2[8 ][ 8: 6],chdata_r2[9 ][ 8: 6],
                     chdata_r2[10 ][ 8: 6],chdata_r2[11 ][ 8: 6],
                     chdata_r2[12 ][ 8: 6],chdata_r2[13 ][ 8: 6],
                     chdata_r2[14 ][ 8: 6],chdata_r2[15][ 8: 6]};
    5'd 3:chdata_o={chdata_r2[0 ][11: 9],chdata_r2[1 ][11: 9],
                     chdata_r2[2 ][11: 9],chdata_r2[3 ][11: 9],
                     chdata_r2[4 ][11: 9],chdata_r2[5 ][11: 9],
                     chdata_r2[6 ][11: 9],chdata_r2[7 ][11: 9],
                     chdata_r2[8 ][11: 9],chdata_r2[9 ][11: 9],
                     chdata_r2[10 ][11: 9],chdata_r2[11 ][11: 9],
                     chdata_r2[12 ][11: 9],chdata_r2[13 ][11: 9],
                     chdata_r2[14 ][11: 9],chdata_r2[15][11: 9]};
    5'd 4:chdata_o={chdata_r2[0 ][14:12],chdata_r2[1 ][14:12],
                     chdata_r2[2 ][14:12],chdata_r2[3 ][14:12],
                     chdata_r2[4 ][14:12],chdata_r2[5 ][14:12],
                     chdata_r2[6 ][14:12],chdata_r2[7 ][14:12],
                     chdata_r2[8 ][14:12],chdata_r2[9 ][14:12],
                     chdata_r2[10 ][14:12],chdata_r2[11 ][14:12],
                     chdata_r2[12 ][14:12],chdata_r2[13 ][14:12],
                     chdata_r2[14 ][14:12],chdata_r2[15][14:12]};
    5'd 5:chdata_o={chdata_r2[0 ][17:15],chdata_r2[1 ][17:15],
                     chdata_r2[2 ][17:15],chdata_r2[3 ][17:15],
                     chdata_r2[4 ][17:15],chdata_r2[5 ][17:15],
                     chdata_r2[6 ][17:15],chdata_r2[7 ][17:15],
                     chdata_r2[8 ][17:15],chdata_r2[9 ][17:15],
                     chdata_r2[10 ][17:15],chdata_r2[11 ][17:15],
                     chdata_r2[12 ][17:15],chdata_r2[13 ][17:15],
                     chdata_r2[14 ][17:15],chdata_r2[15][17:15]};
    5'd 6:chdata_o={chdata_r2[0 ][20:18],chdata_r2[1 ][20:18],
                     chdata_r2[2 ][20:18],chdata_r2[3 ][20:18],
                     chdata_r2[4 ][20:18],chdata_r2[5 ][20:18],
                     chdata_r2[6 ][20:18],chdata_r2[7 ][20:18],
                     chdata_r2[8 ][20:18],chdata_r2[9 ][20:18],
                     chdata_r2[10 ][20:18],chdata_r2[11 ][20:18],
                     chdata_r2[12 ][20:18],chdata_r2[13 ][20:18],
                     chdata_r2[14 ][20:18],chdata_r2[15][20:18]};
    5'd 7:chdata_o={chdata_r2[0 ][23:21],chdata_r2[1 ][23:21],
                     chdata_r2[2 ][23:21],chdata_r2[3 ][23:21],
                     chdata_r2[4 ][23:21],chdata_r2[5 ][23:21],
                     chdata_r2[6 ][23:21],chdata_r2[7 ][23:21],
                     chdata_r2[8 ][23:21],chdata_r2[9 ][23:21],
                     chdata_r2[10 ][23:21],chdata_r2[11 ][23:21],
                     chdata_r2[12 ][23:21],chdata_r2[13 ][23:21],
                     chdata_r2[14 ][23:21],chdata_r2[15][23:21]};
    5'd 8:chdata_o={chdata_r2[0 ][26:24],chdata_r2[1 ][26:24],
                     chdata_r2[2 ][26:24],chdata_r2[3 ][26:24],
                     chdata_r2[4 ][26:24],chdata_r2[5 ][26:24],
                     chdata_r2[6 ][26:24],chdata_r2[7 ][26:24],
                     chdata_r2[8 ][26:24],chdata_r2[9 ][26:24],
                     chdata_r2[10 ][26:24],chdata_r2[11 ][26:24],
                     chdata_r2[12 ][26:24],chdata_r2[13 ][26:24],
                     chdata_r2[14 ][26:24],chdata_r2[15][26:24]};
    5'd 9:chdata_o={chdata_r2[0 ][29:27],chdata_r2[1 ][29:27],
                     chdata_r2[2 ][29:27],chdata_r2[3 ][29:27],
                     chdata_r2[4 ][29:27],chdata_r2[5 ][29:27],
                     chdata_r2[6 ][29:27],chdata_r2[7 ][29:27],
                     chdata_r2[8 ][29:27],chdata_r2[9 ][29:27],
                     chdata_r2[10 ][29:27],chdata_r2[11 ][29:27],
                     chdata_r2[12 ][29:27],chdata_r2[13 ][29:27],
                     chdata_r2[14 ][29:27],chdata_r2[15][29:27]};
    5'd10:chdata_o={chdata_r2[0 ][32:30],chdata_r2[1 ][32:30],
                     chdata_r2[2 ][32:30],chdata_r2[3 ][32:30],
                     chdata_r2[4 ][32:30],chdata_r2[5 ][32:30],
                     chdata_r2[6 ][32:30],chdata_r2[7 ][32:30],
                     chdata_r2[8 ][32:30],chdata_r2[9 ][32:30],
                     chdata_r2[10 ][32:30],chdata_r2[11 ][32:30],
                     chdata_r2[12 ][32:30],chdata_r2[13 ][32:30],
                     chdata_r2[14 ][32:30],chdata_r2[15][32:30]};
    5'd11:chdata_o={chdata_r2[0 ][35:33],chdata_r2[1 ][35:33],
                     chdata_r2[2 ][35:33],chdata_r2[3 ][35:33],
                     chdata_r2[4 ][35:33],chdata_r2[5 ][35:33],
                     chdata_r2[6 ][35:33],chdata_r2[7 ][35:33],
                     chdata_r2[8 ][35:33],chdata_r2[9 ][35:33],
                     chdata_r2[10 ][35:33],chdata_r2[11 ][35:33],
                     chdata_r2[12 ][35:33],chdata_r2[13 ][35:33],
                     chdata_r2[14 ][35:33],chdata_r2[15][35:33]};
    5'd12:chdata_o={chdata_r2[0 ][38:36],chdata_r2[1 ][38:36],
                     chdata_r2[2 ][38:36],chdata_r2[3 ][38:36],
                     chdata_r2[4 ][38:36],chdata_r2[5 ][38:36],
                     chdata_r2[6 ][38:36],chdata_r2[7 ][38:36],
                     chdata_r2[8 ][38:36],chdata_r2[9 ][38:36],
                     chdata_r2[10 ][38:36],chdata_r2[11 ][38:36],
                     chdata_r2[12 ][38:36],chdata_r2[13 ][38:36],
                     chdata_r2[14 ][38:36],chdata_r2[15][38:36]};
    5'd13:chdata_o={chdata_r2[0 ][41:39],chdata_r2[1 ][41:39],
                     chdata_r2[2 ][41:39],chdata_r2[3 ][41:39],
                     chdata_r2[4 ][41:39],chdata_r2[5 ][41:39],
                     chdata_r2[6 ][41:39],chdata_r2[7 ][41:39],
                     chdata_r2[8 ][41:39],chdata_r2[9 ][41:39],
                     chdata_r2[10 ][41:39],chdata_r2[11 ][41:39],
                     chdata_r2[12 ][41:39],chdata_r2[13 ][41:39],
                     chdata_r2[14 ][41:39],chdata_r2[15][41:39]};
    5'd14:chdata_o={chdata_r2[0 ][44:42],chdata_r2[1 ][44:42],
                     chdata_r2[2 ][44:42],chdata_r2[3 ][44:42],
                     chdata_r2[4 ][44:42],chdata_r2[5 ][44:42],
                     chdata_r2[6 ][44:42],chdata_r2[7 ][44:42],
                     chdata_r2[8 ][44:42],chdata_r2[9 ][44:42],
                     chdata_r2[10 ][44:42],chdata_r2[11 ][44:42],
                     chdata_r2[12 ][44:42],chdata_r2[13 ][44:42],
                     chdata_r2[14 ][44:42],chdata_r2[15][44:42]};
    5'd15:chdata_o={chdata_r2[0 ][47:45],chdata_r2[1 ][47:45],
                     chdata_r2[2 ][47:45],chdata_r2[3 ][47:45],
                     chdata_r2[4 ][47:45],chdata_r2[5 ][47:45],
                     chdata_r2[6 ][47:45],chdata_r2[7 ][47:45],
                     chdata_r2[8 ][47:45],chdata_r2[9 ][47:45],
                     chdata_r2[10 ][47:45],chdata_r2[11 ][47:45],
                     chdata_r2[12 ][47:45],chdata_r2[13 ][47:45],
                     chdata_r2[14 ][47:45],chdata_r2[15][47:45]};
    5'd16:chdata_o={chdata_r1[0 ][ 2: 0],chdata_r1[1 ][ 2: 0],
                     chdata_r1[2 ][ 2: 0],chdata_r1[3 ][ 2: 0],
                     chdata_r1[4 ][ 2: 0],chdata_r1[5 ][ 2: 0],
                     chdata_r1[6 ][ 2: 0],chdata_r1[7 ][ 2: 0],
                     chdata_r1[8 ][ 2: 0],chdata_r1[9 ][ 2: 0],
                     chdata_r1[10 ][ 2: 0],chdata_r1[11 ][ 2: 0],
                     chdata_r1[12 ][ 2: 0],chdata_r1[13 ][ 2: 0],
                     chdata_r1[14 ][ 2: 0],chdata_r1[15][ 2: 0]};
    5'd17:chdata_o={chdata_r1[0 ][ 5: 3],chdata_r1[1 ][ 5: 3],
                     chdata_r1[2 ][ 5: 3],chdata_r1[3 ][ 5: 3],
                     chdata_r1[4 ][ 5: 3],chdata_r1[5 ][ 5: 3],
                     chdata_r1[6 ][ 5: 3],chdata_r1[7 ][ 5: 3],
                     chdata_r1[8 ][ 5: 3],chdata_r1[9 ][ 5: 3],
                     chdata_r1[10 ][ 5: 3],chdata_r1[11 ][ 5: 3],
                     chdata_r1[12 ][ 5: 3],chdata_r1[13 ][ 5: 3],
                     chdata_r1[14 ][ 5: 3],chdata_r1[15][ 5: 3]};
    5'd18:chdata_o={chdata_r1[0 ][ 8: 6],chdata_r1[1 ][ 8: 6],
                     chdata_r1[2 ][ 8: 6],chdata_r1[3 ][ 8: 6],
                     chdata_r1[4 ][ 8: 6],chdata_r1[5 ][ 8: 6],
                     chdata_r1[6 ][ 8: 6],chdata_r1[7 ][ 8: 6],
                     chdata_r1[8 ][ 8: 6],chdata_r1[9 ][ 8: 6],
                     chdata_r1[10 ][ 8: 6],chdata_r1[11 ][ 8: 6],
                     chdata_r1[12 ][ 8: 6],chdata_r1[13 ][ 8: 6],
                     chdata_r1[14 ][ 8: 6],chdata_r1[15][ 8: 6]};
    5'd19:chdata_o={chdata_r1[0 ][11: 9],chdata_r1[1 ][11: 9],
                     chdata_r1[2 ][11: 9],chdata_r1[3 ][11: 9],
                     chdata_r1[4 ][11: 9],chdata_r1[5 ][11: 9],
                     chdata_r1[6 ][11: 9],chdata_r1[7 ][11: 9],
                     chdata_r1[8 ][11: 9],chdata_r1[9 ][11: 9],
                     chdata_r1[10 ][11: 9],chdata_r1[11 ][11: 9],
                     chdata_r1[12 ][11: 9],chdata_r1[13 ][11: 9],
                     chdata_r1[14 ][11: 9],chdata_r1[15][11: 9]};
    5'd20:chdata_o={chdata_r1[0 ][14:12],chdata_r1[1 ][14:12],
                     chdata_r1[2 ][14:12],chdata_r1[3 ][14:12],
                     chdata_r1[4 ][14:12],chdata_r1[5 ][14:12],
                     chdata_r1[6 ][14:12],chdata_r1[7 ][14:12],
                     chdata_r1[8 ][14:12],chdata_r1[9 ][14:12],
                     chdata_r1[10 ][14:12],chdata_r1[11 ][14:12],
                     chdata_r1[12 ][14:12],chdata_r1[13 ][14:12],
                     chdata_r1[14 ][14:12],chdata_r1[15][14:12]};
    5'd21:chdata_o={chdata_r1[0 ][17:15],chdata_r1[1 ][17:15],
                     chdata_r1[2 ][17:15],chdata_r1[3 ][17:15],
                     chdata_r1[4 ][17:15],chdata_r1[5 ][17:15],
                     chdata_r1[6 ][17:15],chdata_r1[7 ][17:15],
                     chdata_r1[8 ][17:15],chdata_r1[9 ][17:15],
                     chdata_r1[10 ][17:15],chdata_r1[11 ][17:15],
                     chdata_r1[12 ][17:15],chdata_r1[13 ][17:15],
                     chdata_r1[14 ][17:15],chdata_r1[15][17:15]};
    5'd22:chdata_o={chdata_r1[0 ][20:18],chdata_r1[1 ][20:18],
                     chdata_r1[2 ][20:18],chdata_r1[3 ][20:18],
                     chdata_r1[4 ][20:18],chdata_r1[5 ][20:18],
                     chdata_r1[6 ][20:18],chdata_r1[7 ][20:18],
                     chdata_r1[8 ][20:18],chdata_r1[9 ][20:18],
                     chdata_r1[10 ][20:18],chdata_r1[11 ][20:18],
                     chdata_r1[12 ][20:18],chdata_r1[13 ][20:18],
                     chdata_r1[14 ][20:18],chdata_r1[15][20:18]};
    5'd23:chdata_o={chdata_r1[0 ][23:21],chdata_r1[1 ][23:21],
                     chdata_r1[2 ][23:21],chdata_r1[3 ][23:21],
                     chdata_r1[4 ][23:21],chdata_r1[5 ][23:21],
                     chdata_r1[6 ][23:21],chdata_r1[7 ][23:21],
                     chdata_r1[8 ][23:21],chdata_r1[9 ][23:21],
                     chdata_r1[10 ][23:21],chdata_r1[11 ][23:21],
                     chdata_r1[12 ][23:21],chdata_r1[13 ][23:21],
                     chdata_r1[14 ][23:21],chdata_r1[15][23:21]};
    5'd24:chdata_o={chdata_r1[0 ][26:24],chdata_r1[1 ][26:24],
                     chdata_r1[2 ][26:24],chdata_r1[3 ][26:24],
                     chdata_r1[4 ][26:24],chdata_r1[5 ][26:24],
                     chdata_r1[6 ][26:24],chdata_r1[7 ][26:24],
                     chdata_r1[8 ][26:24],chdata_r1[9 ][26:24],
                     chdata_r1[10 ][26:24],chdata_r1[11 ][26:24],
                     chdata_r1[12 ][26:24],chdata_r1[13 ][26:24],
                     chdata_r1[14 ][26:24],chdata_r1[15][26:24]};
    5'd25:chdata_o={chdata_r1[0 ][29:27],chdata_r1[1 ][29:27],
                     chdata_r1[2 ][29:27],chdata_r1[3 ][29:27],
                     chdata_r1[4 ][29:27],chdata_r1[5 ][29:27],
                     chdata_r1[6 ][29:27],chdata_r1[7 ][29:27],
                     chdata_r1[8 ][29:27],chdata_r1[9 ][29:27],
                     chdata_r1[10 ][29:27],chdata_r1[11 ][29:27],
                     chdata_r1[12 ][29:27],chdata_r1[13 ][29:27],
                     chdata_r1[14 ][29:27],chdata_r1[15][29:27]};
    5'd26:chdata_o={chdata_r1[0 ][32:30],chdata_r1[1 ][32:30],
                     chdata_r1[2 ][32:30],chdata_r1[3 ][32:30],
                     chdata_r1[4 ][32:30],chdata_r1[5 ][32:30],
                     chdata_r1[6 ][32:30],chdata_r1[7 ][32:30],
                     chdata_r1[8 ][32:30],chdata_r1[9 ][32:30],
                     chdata_r1[10 ][32:30],chdata_r1[11 ][32:30],
                     chdata_r1[12 ][32:30],chdata_r1[13 ][32:30],
                     chdata_r1[14 ][32:30],chdata_r1[15][32:30]};
    5'd27:chdata_o={chdata_r1[0 ][35:33],chdata_r1[1 ][35:33],
                     chdata_r1[2 ][35:33],chdata_r1[3 ][35:33],
                     chdata_r1[4 ][35:33],chdata_r1[5 ][35:33],
                     chdata_r1[6 ][35:33],chdata_r1[7 ][35:33],
                     chdata_r1[8 ][35:33],chdata_r1[9 ][35:33],
                     chdata_r1[10 ][35:33],chdata_r1[11 ][35:33],
                     chdata_r1[12 ][35:33],chdata_r1[13 ][35:33],
                     chdata_r1[14 ][35:33],chdata_r1[15][35:33]};
    5'd28:chdata_o={chdata_r1[0 ][38:36],chdata_r1[1 ][38:36],
                     chdata_r1[2 ][38:36],chdata_r1[3 ][38:36],
                     chdata_r1[4 ][38:36],chdata_r1[5 ][38:36],
                     chdata_r1[6 ][38:36],chdata_r1[7 ][38:36],
                     chdata_r1[8 ][38:36],chdata_r1[9 ][38:36],
                     chdata_r1[10 ][38:36],chdata_r1[11 ][38:36],
                     chdata_r1[12 ][38:36],chdata_r1[13 ][38:36],
                     chdata_r1[14 ][38:36],chdata_r1[15][38:36]};
    5'd29:chdata_o={chdata_r1[0 ][41:39],chdata_r1[1 ][41:39],
                     chdata_r1[2 ][41:39],chdata_r1[3 ][41:39],
                     chdata_r1[4 ][41:39],chdata_r1[5 ][41:39],
                     chdata_r1[6 ][41:39],chdata_r1[7 ][41:39],
                     chdata_r1[8 ][41:39],chdata_r1[9 ][41:39],
                     chdata_r1[10 ][41:39],chdata_r1[11 ][41:39],
                     chdata_r1[12 ][41:39],chdata_r1[13 ][41:39],
                     chdata_r1[14 ][41:39],chdata_r1[15][41:39]};
    5'd30:chdata_o={chdata_r1[0 ][44:42],chdata_r1[1 ][44:42],
                     chdata_r1[2 ][44:42],chdata_r1[3 ][44:42],
                     chdata_r1[4 ][44:42],chdata_r1[5 ][44:42],
                     chdata_r1[6 ][44:42],chdata_r1[7 ][44:42],
                     chdata_r1[8 ][44:42],chdata_r1[9 ][44:42],
                     chdata_r1[10 ][44:42],chdata_r1[11 ][44:42],
                     chdata_r1[12 ][44:42],chdata_r1[13 ][44:42],
                     chdata_r1[14 ][44:42],chdata_r1[15][44:42]};
    5'd31:chdata_o={chdata_r1[0 ][47:45],chdata_r1[1 ][47:45],
                     chdata_r1[2 ][47:45],chdata_r1[3 ][47:45],
                     chdata_r1[4 ][47:45],chdata_r1[5 ][47:45],
                     chdata_r1[6 ][47:45],chdata_r1[7 ][47:45],
                     chdata_r1[8 ][47:45],chdata_r1[9 ][47:45],
                     chdata_r1[10 ][47:45],chdata_r1[11 ][47:45],
                     chdata_r1[12 ][47:45],chdata_r1[13 ][47:45],
                     chdata_r1[14 ][47:45],chdata_r1[15][47:45]};
    default: chdata_o=0;
  endcase
end
always @(negedge RESET_N or posedge CLK)
if (~RESET_N)
begin
  counter <=0;
  memid   <=0;
  memgroup<=0;
  section_ch<=0;
end
else
begin
  counter<=((~data_wrsa & ~data_wrsb)| (counter==5'd31))?
            5'd0:counter+5'd1;
  if(load_data_en)
  begin
    section_ch  <=(counter==5'd15 | counter==5'd31)?section_ch+2'd1:section_ch;
  if(counter==5'd15 | counter==5'd31)
    memid<=(memid==3'd7)? 3'd0 :
           (~data_wrsa & ~data_wrsb)? 3'd0 : memid+3'd1;
  if(section_ch==2'd3 & memid==3'd7 & (counter==5'd15 | counter==5'd31))
    memgroup<=(memgroup==3'd4)?
               3'd5 : memgroup+3'd1;
  end
  else
  begin
    memid     <=0;
    memgroup  <=0;
    section_ch<=0;
  end
end
integer i;
always @(negedge RESET_N or posedge CLK)
if (~RESET_N)
begin
  for (i=0; i<=15; i=i+1)  chdata_r1[i ]<=0;
  for (i=0; i<=15; i=i+1)  chdata_r2[i ]<=0;
end
else
begin
  case(counter)
    5'd0:chdata_r1 [0] <=chdata_w;
    5'd1:chdata_r1 [1] <=chdata_w;
    5'd2:chdata_r1 [2] <=chdata_w;
    5'd3:chdata_r1 [3] <=chdata_w;
    5'd4:chdata_r1 [4] <=chdata_w;
    5'd5:chdata_r1 [5] <=chdata_w;
    5'd6:chdata_r1 [6] <=chdata_w;
    5'd7:chdata_r1 [7] <=chdata_w;
    5'd8:chdata_r1 [8] <=chdata_w;
    5'd9:chdata_r1 [9] <=chdata_w;
    5'd10:chdata_r1[10]<=chdata_w;
    5'd11:chdata_r1[11]<=chdata_w;
    5'd12:chdata_r1[12]<=chdata_w;
    5'd13:chdata_r1[13]<=chdata_w;
    5'd14:chdata_r1[14]<=chdata_w;
    5'd15:chdata_r1[15]<=chdata_w;
    5'd16:chdata_r2[0] <=chdata_w;
    5'd17:chdata_r2[1] <=chdata_w;
    5'd18:chdata_r2[2] <=chdata_w;
    5'd19:chdata_r2[3] <=chdata_w;
    5'd20:chdata_r2[4] <=chdata_w;
    5'd21:chdata_r2[5] <=chdata_w;
    5'd22:chdata_r2[6] <=chdata_w;
    5'd23:chdata_r2[7] <=chdata_w;
    5'd24:chdata_r2[8] <=chdata_w;
    5'd25:chdata_r2[9] <=chdata_w;
    5'd26:chdata_r2[10]<=chdata_w;
    5'd27:chdata_r2[11]<=chdata_w;
    5'd28:chdata_r2[12]<=chdata_w;
    5'd29:chdata_r2[13]<=chdata_w;
    5'd30:chdata_r2[14]<=chdata_w;
    5'd31:chdata_r2[15]<=chdata_w;
  endcase
end
endmodule

module  invrotatreg(
                 CLK,RESET_N,
                 hb_en,start_ldpc,
                 data_wrsa,data_wrsb,
                 hbout,
                 hbout_o);

input CLK,RESET_N,hb_en,start_ldpc,
      data_wrsa,data_wrsb;
input [15:0] hbout;
output [15:0] hbout_o;
reg [4:0] counter;
reg [15:0] hbout_r1,hbout_r2,hbout_r3,hbout_r4,
           hbout_r5,hbout_r6,hbout_r7,hbout_r8,
                 hbout_r9,hbout_r10,hbout_r11,hbout_r12,
                 hbout_r13,hbout_r14,hbout_r15,hbout_r16,
                 hbout_r17,hbout_r18,hbout_r19,hbout_r20,
                 hbout_r21,hbout_r22,hbout_r23,hbout_r24,
                 hbout_r25,hbout_r26,hbout_r27,hbout_r28,
                 hbout_r29,hbout_r30,hbout_r31,hbout_r32;
reg [15:0] hbout_o;
reg [1:0] section_hb;

always @(*)
begin
  case(counter)
    5'd 1:hbout_o={hbout_r32[0 ],hbout_r31[0 ],hbout_r30[0 ],hbout_r29[0 ],
                   hbout_r28[0 ],hbout_r27[0 ],hbout_r26[0 ],hbout_r25[0 ],
                   hbout_r24[0 ],hbout_r23[0 ],hbout_r22[ 0],hbout_r21[0 ],
                   hbout_r20[0 ],hbout_r19[0 ],hbout_r18[0 ],hbout_r17[0 ]};
    5'd 2:hbout_o={
                   hbout_r32[1],hbout_r31[1],hbout_r30[1],hbout_r29[1],
                   hbout_r28[1],hbout_r27[1],hbout_r26[1],hbout_r25[1],
                   hbout_r24[1],hbout_r23[1],hbout_r22[1],hbout_r21[1],
                   hbout_r20[1],hbout_r19[1],hbout_r18[1],hbout_r17[1]};
    5'd 3:hbout_o={
                   hbout_r32[2],hbout_r31[2],hbout_r30[2],hbout_r29[2],
                   hbout_r28[2],hbout_r27[2],hbout_r26[2],hbout_r25[2],
                   hbout_r24[2],hbout_r23[2],hbout_r22[2],hbout_r21[2],
                   hbout_r20[2],hbout_r19[2],hbout_r18[2],hbout_r17[2]};
    5'd 4:hbout_o={
                   hbout_r32[3],hbout_r31[3],hbout_r30[3],hbout_r29[3],
                   hbout_r28[3],hbout_r27[3],hbout_r26[3],hbout_r25[3],
                   hbout_r24[3],hbout_r23[3],hbout_r22[3],hbout_r21[3],
                   hbout_r20[3],hbout_r19[3],hbout_r18[3],hbout_r17[3]};
    5'd 5:hbout_o={
                   hbout_r32[4],hbout_r31[4],hbout_r30[4],hbout_r29[4],
                   hbout_r28[4],hbout_r27[4],hbout_r26[4],hbout_r25[4],
                   hbout_r24[4],hbout_r23[4],hbout_r22[4],hbout_r21[4],
                   hbout_r20[4],hbout_r19[4],hbout_r18[4],hbout_r17[4]};
    5'd 6:hbout_o={
                   hbout_r32[5],hbout_r31[5],hbout_r30[5],hbout_r29[5],
                   hbout_r28[5],hbout_r27[5],hbout_r26[5],hbout_r25[5],
                   hbout_r24[5],hbout_r23[5],hbout_r22[5],hbout_r21[5],
                   hbout_r20[5],hbout_r19[5],hbout_r18[5],hbout_r17[5]};
    5'd 7:hbout_o={
                   hbout_r32[6],hbout_r31[6],hbout_r30[6],hbout_r29[6],
                   hbout_r28[6],hbout_r27[6],hbout_r26[6],hbout_r25[6],
                   hbout_r24[6],hbout_r23[6],hbout_r22[6],hbout_r21[6],
                   hbout_r20[6],hbout_r19[6],hbout_r18[6],hbout_r17[6]};
    5'd 8:hbout_o={
                   hbout_r32[7],hbout_r31[7],hbout_r30[7],hbout_r29[7],
                   hbout_r28[7],hbout_r27[7],hbout_r26[7],hbout_r25[7],
                   hbout_r24[7],hbout_r23[7],hbout_r22[7],hbout_r21[7],
                   hbout_r20[7],hbout_r19[7],hbout_r18[7],hbout_r17[7]};
    5'd 9:hbout_o={
                   hbout_r32[8],hbout_r31[8],hbout_r30[8],hbout_r29[8],
                   hbout_r28[8],hbout_r27[8],hbout_r26[8],hbout_r25[8],
                   hbout_r24[8],hbout_r23[8],hbout_r22[8],hbout_r21[8],
                   hbout_r20[8],hbout_r19[8],hbout_r18[8],hbout_r17[8]};
    5'd10:hbout_o={
                   hbout_r32[9],hbout_r31[9],hbout_r30[9],hbout_r29[9],
                   hbout_r28[9],hbout_r27[9],hbout_r26[9],hbout_r25[9],
                   hbout_r24[9],hbout_r23[9],hbout_r22[9],hbout_r21[9],
                   hbout_r20[9],hbout_r19[9],hbout_r18[9],hbout_r17[9]};
    5'd11:hbout_o={
                   hbout_r32[10],hbout_r31[10],hbout_r30[10],hbout_r29[10],
                   hbout_r28[10],hbout_r27[10],hbout_r26[10],hbout_r25[10],
                   hbout_r24[10],hbout_r23[10],hbout_r22[10],hbout_r21[10],
                   hbout_r20[10],hbout_r19[10],hbout_r18[10],hbout_r17[10]};
    5'd12:hbout_o={
                   hbout_r32[11],hbout_r31[11],hbout_r30[11],hbout_r29[11],
                   hbout_r28[11],hbout_r27[11],hbout_r26[11],hbout_r25[11],
                   hbout_r24[11],hbout_r23[11],hbout_r22[11],hbout_r21[11],
                   hbout_r20[11],hbout_r19[11],hbout_r18[11],hbout_r17[11]};
    5'd13:hbout_o={
                   hbout_r32[12],hbout_r31[12],hbout_r30[12],hbout_r29[12],
                   hbout_r28[12],hbout_r27[12],hbout_r26[12],hbout_r25[12],
                   hbout_r24[12],hbout_r23[12],hbout_r22[12],hbout_r21[12],
                   hbout_r20[12],hbout_r19[12],hbout_r18[12],hbout_r17[12]};
    5'd14:hbout_o={
                   hbout_r32[13],hbout_r31[13],hbout_r30[13],hbout_r29[13],
                   hbout_r28[13],hbout_r27[13],hbout_r26[13],hbout_r25[13],
                   hbout_r24[13],hbout_r23[13],hbout_r22[13],hbout_r21[13],
                   hbout_r20[13],hbout_r19[13],hbout_r18[13],hbout_r17[13]};
    5'd15:hbout_o={
                   hbout_r32[14],hbout_r31[14],hbout_r30[14],hbout_r29[14],
                   hbout_r28[14],hbout_r27[14],hbout_r26[14],hbout_r25[14],
                   hbout_r24[14],hbout_r23[14],hbout_r22[14],hbout_r21[14],
                   hbout_r20[14],hbout_r19[14],hbout_r18[14],hbout_r17[14]};
    5'd16:hbout_o={
                   hbout_r32[15],hbout_r31[15],hbout_r30[15],hbout_r29[15],
                   hbout_r28[15],hbout_r27[15],hbout_r26[15],hbout_r25[15],
                   hbout_r24[15],hbout_r23[15],hbout_r22[15],hbout_r21[15],
                   hbout_r20[15],hbout_r19[15],hbout_r18[15],hbout_r17[15]};
    5'd17:hbout_o={
                   hbout_r16[0 ],hbout_r15[0 ],hbout_r14[0 ],hbout_r13[0 ],
                   hbout_r12[0 ],hbout_r11[0 ],hbout_r10[0 ],hbout_r9 [0 ],
                   hbout_r8 [0 ],hbout_r7 [0 ],hbout_r6 [0 ],hbout_r5 [0 ],
                   hbout_r4 [0 ],hbout_r3 [0 ],hbout_r2 [0 ],hbout_r1 [0 ]};
    5'd18:hbout_o={
                   hbout_r16[1 ],hbout_r15[1 ],hbout_r14[1 ],hbout_r13[1 ],
                   hbout_r12[1 ],hbout_r11[1 ],hbout_r10[1 ],hbout_r9 [1 ],
                   hbout_r8 [1 ],hbout_r7 [1 ],hbout_r6 [1 ],hbout_r5 [1 ],
                   hbout_r4 [1 ],hbout_r3 [1 ],hbout_r2 [1 ],hbout_r1 [1 ]};
    5'd19:hbout_o={
                   hbout_r16[2 ],hbout_r15[2 ],hbout_r14[2 ],hbout_r13[2 ],
                   hbout_r12[2 ],hbout_r11[2 ],hbout_r10[2 ],hbout_r9 [2 ],
                   hbout_r8 [2 ],hbout_r7 [2 ],hbout_r6 [2 ],hbout_r5 [2 ],
                   hbout_r4 [2 ],hbout_r3 [2 ],hbout_r2 [2 ],hbout_r1 [2 ]};
    5'd20:hbout_o={
                   hbout_r16[3 ],hbout_r15[3 ],hbout_r14[3 ],hbout_r13[3 ],
                   hbout_r12[3 ],hbout_r11[3 ],hbout_r10[3 ],hbout_r9 [3 ],
                   hbout_r8 [3 ],hbout_r7 [3 ],hbout_r6 [3 ],hbout_r5 [3 ],
                   hbout_r4 [3 ],hbout_r3 [3 ],hbout_r2 [3 ],hbout_r1 [3 ]};
    5'd21:hbout_o={
                   hbout_r16[4 ],hbout_r15[4 ],hbout_r14[4 ],hbout_r13[4 ],
                   hbout_r12[4 ],hbout_r11[4 ],hbout_r10[4 ],hbout_r9 [4 ],
                   hbout_r8 [4 ],hbout_r7 [4 ],hbout_r6 [4 ],hbout_r5 [4 ],
                   hbout_r4 [4 ],hbout_r3 [4 ],hbout_r2 [4 ],hbout_r1 [4 ]};
    5'd22:hbout_o={
                   hbout_r16[5 ],hbout_r15[5 ],hbout_r14[5],hbout_r13[5],
                   hbout_r12[5 ],hbout_r11[5 ],hbout_r10[5],hbout_r9 [5],
                   hbout_r8 [5 ],hbout_r7 [5 ],hbout_r6 [5],hbout_r5 [5],
                   hbout_r4 [5 ],hbout_r3 [5 ],hbout_r2 [5],hbout_r1 [5]};
    5'd23:hbout_o={
                   hbout_r16[6 ],hbout_r15[6 ],hbout_r14[6 ],hbout_r13[6],
                   hbout_r12[6 ],hbout_r11[6 ],hbout_r10[6 ],hbout_r9 [6],
                   hbout_r8 [6 ],hbout_r7 [6 ],hbout_r6 [6 ],hbout_r5 [6],
                   hbout_r4 [6 ],hbout_r3 [6 ],hbout_r2 [6 ],hbout_r1 [6]};
    5'd24:hbout_o={
                   hbout_r16[7],hbout_r15[7],hbout_r14[7],hbout_r13[7],
                   hbout_r12[7],hbout_r11[7],hbout_r10[7],hbout_r9 [7],
                   hbout_r8 [7],hbout_r7 [7],hbout_r6 [7],hbout_r5 [7],
                   hbout_r4 [7],hbout_r3 [7],hbout_r2 [7],hbout_r1 [7]};
    5'd25:hbout_o={
                   hbout_r16[8],hbout_r15[8],hbout_r14[8],hbout_r13[8],
                   hbout_r12[8],hbout_r11[8],hbout_r10[8],hbout_r9 [8],
                   hbout_r8 [8],hbout_r7 [8],hbout_r6 [8],hbout_r5 [8],
                   hbout_r4 [8],hbout_r3 [8],hbout_r2 [8],hbout_r1 [8]};
    5'd26:hbout_o={
                   hbout_r16[9],hbout_r15[9],hbout_r14[9],hbout_r13[9],
                   hbout_r12[9],hbout_r11[9],hbout_r10[9],hbout_r9 [9],
                   hbout_r8 [9],hbout_r7 [9],hbout_r6 [9],hbout_r5 [9],
                   hbout_r4 [9],hbout_r3 [9],hbout_r2 [9],hbout_r1 [9]};
    5'd27:hbout_o={
                   hbout_r16[10],hbout_r15[10],hbout_r14[10],hbout_r13[10],
                   hbout_r12[10],hbout_r11[10],hbout_r10[10],hbout_r9 [10],
                   hbout_r8 [10],hbout_r7 [10],hbout_r6 [10],hbout_r5 [10],
                   hbout_r4 [10],hbout_r3 [10],hbout_r2 [10],hbout_r1 [10]};
    5'd28:hbout_o={
                   hbout_r16[11],hbout_r15[11],hbout_r14[11],hbout_r13[11],
                   hbout_r12[11],hbout_r11[11],hbout_r10[11],hbout_r9 [11],
                   hbout_r8 [11],hbout_r7 [11],hbout_r6 [11],hbout_r5 [11],
                   hbout_r4 [11],hbout_r3 [11],hbout_r2 [11],hbout_r1 [11]};
    5'd29:hbout_o={
                   hbout_r16[12],hbout_r15[12],hbout_r14[12],hbout_r13[12],
                   hbout_r12[12],hbout_r11[12],hbout_r10[12],hbout_r9 [12],
                   hbout_r8 [12],hbout_r7 [12],hbout_r6 [12],hbout_r5 [12],
                   hbout_r4 [12],hbout_r3 [12],hbout_r2 [12],hbout_r1 [12]};
    5'd30:hbout_o={
                   hbout_r16[13],hbout_r15[13],hbout_r14[13],hbout_r13[13],
                   hbout_r12[13],hbout_r11[13],hbout_r10[13],hbout_r9 [13],
                   hbout_r8 [13],hbout_r7 [13],hbout_r6 [13],hbout_r5 [13],
                   hbout_r4 [13],hbout_r3 [13],hbout_r2 [13],hbout_r1 [13]};
    5'd31:hbout_o={
                   hbout_r16[14],hbout_r15[14],hbout_r14[14],hbout_r13[14],
                   hbout_r12[14],hbout_r11[14],hbout_r10[14],hbout_r9 [14],
                   hbout_r8 [14],hbout_r7 [14],hbout_r6 [14],hbout_r5 [14],
                   hbout_r4 [14],hbout_r3 [14],hbout_r2 [14],hbout_r1 [14]};
    5'd0:hbout_o={hbout_r16[15],hbout_r15[15],hbout_r14[15],hbout_r13[15],
                   hbout_r12[15],hbout_r11[15],hbout_r10[15],hbout_r9 [15],
                   hbout_r8 [15],hbout_r7 [15],hbout_r6 [15],hbout_r5 [15],
                   hbout_r4 [15],hbout_r3 [15],hbout_r2 [15],hbout_r1 [15]};
    default: hbout_o=0;
  endcase
end
always @(negedge RESET_N or posedge CLK)
if (~RESET_N)
begin
  counter <=0;
end
else
begin
  counter<=(hb_en)?((counter==5'd31)?
            5'd0:counter+5'd1):5'd0;
end

always @(negedge RESET_N or posedge CLK)
if (~RESET_N)
begin
   hbout_r1 <=0;
   hbout_r2 <=0;
   hbout_r3 <=0;
   hbout_r4 <=0;
   hbout_r5 <=0;
   hbout_r6 <=0;
   hbout_r7 <=0;
   hbout_r8 <=0;
   hbout_r9 <=0;
   hbout_r10<=0;
   hbout_r11<=0;
   hbout_r12<=0;
   hbout_r13<=0;
   hbout_r14<=0;
   hbout_r15<=0;
   hbout_r16<=0;
   hbout_r17<=0;
   hbout_r18<=0;
   hbout_r19<=0;
   hbout_r20<=0;
   hbout_r21<=0;
   hbout_r22<=0;
   hbout_r23<=0;
   hbout_r24<=0;
   hbout_r25<=0;
   hbout_r26<=0;
   hbout_r27<=0;
   hbout_r28<=0;
   hbout_r29<=0;
   hbout_r30<=0;
   hbout_r31<=0;
   hbout_r32<=0;
end
else
begin
  if(hb_en)
  begin
  case(counter)
    5'd 1:hbout_r1 <=hbout;
    5'd 2:hbout_r2 <=hbout;
    5'd 3:hbout_r3 <=hbout;
    5'd 4:hbout_r4 <=hbout;
    5'd 5:hbout_r5 <=hbout;
    5'd 6:hbout_r6 <=hbout;
    5'd 7:hbout_r7 <=hbout;
    5'd 8:hbout_r8 <=hbout;
    5'd 9:hbout_r9 <=hbout;
    5'd10:hbout_r10<=hbout;
    5'd11:hbout_r11<=hbout;
    5'd12:hbout_r12<=hbout;
    5'd13:hbout_r13<=hbout;
    5'd14:hbout_r14<=hbout;
    5'd15:hbout_r15<=hbout;
    5'd16:hbout_r16<=hbout;
    5'd17:hbout_r17<=hbout;
    5'd18:hbout_r18<=hbout;
    5'd19:hbout_r19<=hbout;
    5'd20:hbout_r20<=hbout;
    5'd21:hbout_r21<=hbout;
    5'd22:hbout_r22<=hbout;
    5'd23:hbout_r23<=hbout;
    5'd24:hbout_r24<=hbout;
    5'd25:hbout_r25<=hbout;
    5'd26:hbout_r26<=hbout;
    5'd27:hbout_r27<=hbout;
    5'd28:hbout_r28<=hbout;
    5'd29:hbout_r29<=hbout;
    5'd30:hbout_r30<=hbout;
    5'd31:hbout_r31<=hbout;
    5'd0 :hbout_r32<=hbout;
    default:
    begin
      hbout_r1<=0;
      hbout_r2<=0;
      hbout_r3<=0;
      hbout_r4<=0;
      hbout_r5<=0;
      hbout_r6<=0;
      hbout_r7<=0;
      hbout_r8<=0;
      hbout_r9<=0;
      hbout_r10<=0;
      hbout_r11<=0;
      hbout_r12<=0;
      hbout_r13<=0;
      hbout_r14<=0;
      hbout_r15<=0;
      hbout_r16<=0;
      hbout_r17<=0;
      hbout_r18<=0;
      hbout_r19<=0;
      hbout_r20<=0;
      hbout_r21<=0;
      hbout_r22<=0;
      hbout_r23<=0;
      hbout_r24<=0;
      hbout_r25<=0;
      hbout_r26<=0;
      hbout_r27<=0;
      hbout_r28<=0;
      hbout_r29<=0;
      hbout_r30<=0;
      hbout_r31<=0;
      hbout_r32<=0;
    end
  endcase
 end
end
endmodule

module invpermutator1(
                   section,layer_i,
                   mtv1,mtv2,
                   ctm1_i,ctm2_i,
                   mtv1_w,mtv2_w,
                   sumdata1,sumdata2,sumdata1_w,sumdata2_w,
                   rotat_en,
                   ctm1,ctm2);

input [1:0] layer_i,section;
input [79:0] mtv1,mtv2;
input [47:0] ctm1_i,ctm2_i;
input [79:0] sumdata1,sumdata2;
input [7:0]rotat_en;
output [47:0] ctm1,ctm2;
output [79:0] mtv1_w,mtv2_w;
output [79:0] sumdata1_w,sumdata2_w;

//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//            2st row block   3st row block    4st row block
// shift Ext number  0           0             0
// shift Ext number  3           13            14
// shift Ext number  11          7             12
// shift Ext number  9           8             13
// shift Ext number  1           6             3
// shift Ext number  6           3             15
// shift Ext number  12          13            6
// shift Ext number  3           9             15
wire [47:0]
  ctm1_w=ctm1_i,

  ctm2_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[1])?{ctm1_i[11:0],ctm1_i[47:12]} : {ctm1_i[8:0],ctm1_i[47:9]} :
         (layer_i==2'b10)?(rotat_en[1])?{ctm1_i[41:0],ctm1_i[47:42]} : {ctm1_i[38:0],ctm1_i[47:39]} :
                          (rotat_en[1])?{ctm1_i[44:0],ctm1_i[47:45]} : {ctm1_i[41:0],ctm1_i[47:42]} ,
  ctm3_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[2])?{ctm1_i[35:0],ctm1_i[47:36]} : {ctm1_i[32:0],ctm1_i[47:33]} :
         (layer_i==2'b10)?(rotat_en[2])?{ctm1_i[23:0],ctm1_i[47:24]} : {ctm1_i[20:0],ctm1_i[47:21]} :
                          (rotat_en[2])?{ctm1_i[38:0],ctm1_i[47:39]} : {ctm1_i[35:0],ctm1_i[47:36]} ,
  ctm4_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[3])?{ctm1_i[29:0],ctm1_i[47:30]} : {ctm1_i[26:0],ctm1_i[47:27]} :
         (layer_i==2'b10)?(rotat_en[3])?{ctm1_i[26:0],ctm1_i[47:27]} : {ctm1_i[23:0],ctm1_i[47:24]} :
                          (rotat_en[3])?{ctm1_i[41:0],ctm1_i[47:42]} : {ctm1_i[38:0],ctm1_i[47:39]} ,
  ctm5_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[4])?{ctm2_i[5:0],ctm2_i[47:6]} : {ctm2_i[2:0],ctm2_i[47:3]} :
         (layer_i==2'b10)?(rotat_en[4])?{ctm2_i[20:0],ctm2_i[47:21]} : {ctm2_i[17:0],ctm2_i[47:18]} :
                          (rotat_en[4])?{ctm2_i[11:0],ctm2_i[47:12]} : {ctm2_i[8:0],ctm2_i[47:9]} ,
  ctm6_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[5])?{ctm2_i[20:0],ctm2_i[47:21]} : {ctm2_i[17:0],ctm2_i[47:18]} :
         (layer_i==2'b10)?(rotat_en[5])?{ctm2_i[11:0],ctm2_i[47:12]} : {ctm2_i[8:0],ctm2_i[47:9]} :
                          (rotat_en[5])? ctm2_i : {ctm2_i[44:0],ctm2_i[47:45]} ,
  ctm7_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[6])?{ctm2_i[38:0],ctm2_i[47:39]} : {ctm2_i[35:0],ctm2_i[47:36]} :
         (layer_i==2'b10)?(rotat_en[6])?{ctm2_i[41:0],ctm2_i[47:42]} : {ctm2_i[38:0],ctm2_i[47:39]} :
                          (rotat_en[6])?{ctm2_i[20:0],ctm2_i[47:21]} : {ctm2_i[17:0],ctm2_i[47:18]} ,
  ctm8_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[7])?{ctm2_i[11:0],ctm2_i[47:12]} : {ctm2_i[8:0],ctm2_i[47:9]} :
         (layer_i==2'b10)?(rotat_en[7])?{ctm2_i[29:0],ctm2_i[47:30]} : {ctm2_i[26:0],ctm2_i[47:27]} :
                          (rotat_en[7])? ctm2_i : {ctm2_i[44:0],ctm2_i[47:45]} ;
wire [47:0]
     ctm1=(section==2'b00)?ctm1_w:
          (section==2'b01)?ctm2_w:
          (section==2'b10)?ctm3_w:
                           ctm4_w,
     ctm2=(section==2'b00)?ctm5_w:
          (section==2'b01)?ctm6_w:
          (section==2'b10)?ctm7_w:
                           ctm8_w;
 //            2st row block   3st row block    4st row block
// shift Ext number  0           0             0
// shift Ext number  3           13            14
// shift Ext number  11          7             12
// shift Ext number  9           8             13
// shift Ext number  1           6             3
// shift Ext number  6           3             15
// shift Ext number  12          13            6
// shift Ext number  3           9             15
wire [79:0]         // error
  mtv1w = mtv1,
  mtv2w = (layer_i==2'b00)? mtv1:
          (layer_i==2'b01)? (rotat_en[1])?{mtv1[59:0],mtv1[79:60]} : {mtv1[64:0],mtv1[79:65]}:
          (layer_i==2'b10)? (rotat_en[1])?{mtv1[9:0],mtv1[79:10]} : {mtv1[14:0],mtv1[79:15]} :
                            (rotat_en[1])?{mtv1[4:0],mtv1[79:5]} : {mtv1[9:0],mtv1[79:10]}   ,
  mtv3w = (layer_i==2'b00)? mtv1:
          (layer_i==2'b01)? (rotat_en[2])?{mtv1[19:0],mtv1[79:20]} : {mtv1[24:0],mtv1[79:25]}:
          (layer_i==2'b10)? (rotat_en[2])?{mtv1[39:0],mtv1[79:40]} : {mtv1[44:0],mtv1[79:45]}:
                            (rotat_en[2])?{mtv1[14:0],mtv1[79:15]} : {mtv1[19:0],mtv1[79:20]},
  mtv4w = (layer_i==2'b00)? mtv1:
          (layer_i==2'b01)? (rotat_en[3])?{mtv1[29:0],mtv1[79:30]} : {mtv1[34:0],mtv1[79:35]}:
          (layer_i==2'b10)? (rotat_en[3])?{mtv1[34:0],mtv1[79:35]} : {mtv1[39:0],mtv1[79:40]}:
                            (rotat_en[3])?{mtv1[9:0],mtv1[79:10]} : {mtv1[14:0],mtv1[79:15]} ,
  mtv5w = (layer_i==2'b00)? mtv2:
          (layer_i==2'b01)? (rotat_en[4])?{mtv2[69:0],mtv2[79:70]} : {mtv2[74:0],mtv2[79:75]}:
          (layer_i==2'b10)? (rotat_en[4])?{mtv2[44:0],mtv2[79:45]} : {mtv2[49:0],mtv2[79:50]}:
                            (rotat_en[4])?{mtv2[59:0],mtv2[79:60]} : {mtv2[64:0],mtv2[79:65]},
  mtv6w = (layer_i==2'b00)? mtv2:
          (layer_i==2'b01)? (rotat_en[5])?{mtv2[44:0],mtv2[79:45]} : {mtv2[49:0],mtv2[79:50]}:
          (layer_i==2'b10)? (rotat_en[5])?{mtv2[59:0],mtv2[79:60]} : {mtv2[64:0],mtv2[79:65]}:
                            (rotat_en[5])? mtv2  : {mtv2[4:0],mtv2[79:5]}                        ,
  mtv7w = (layer_i==2'b00)? mtv2:
          (layer_i==2'b01)? (rotat_en[6])?{mtv2[14:0],mtv2[79:15]} : {mtv2[19:0],mtv2[79:20]}:
          (layer_i==2'b10)? (rotat_en[6])?{mtv2[9:0],mtv2[79:10]} : {mtv2[14:0],mtv2[79:15]} :
                            (rotat_en[6])?{mtv2[44:0],mtv2[79:45]} : {mtv2[49:0],mtv2[79:50]},
  mtv8w = (layer_i==2'b00)? mtv2:
          (layer_i==2'b01)? (rotat_en[7])?{mtv2[59:0],mtv2[79:60]} : {mtv2[64:0],mtv2[79:65]}:
          (layer_i==2'b10)? (rotat_en[7])?{mtv2[29:0],mtv2[79:30]} : {mtv2[34:0],mtv2[79:35]}:
                            (rotat_en[7])? mtv2 : {mtv2[4:0],mtv2[79:5]}                         ;

wire [79:0]
  mtv1_w=(section==2'b00)? mtv1w:
         (section==2'b01)? mtv2w:
         (section==2'b10)? mtv3w:
                           mtv4w,
  mtv2_w=(section==2'b00)? mtv5w:
         (section==2'b01)? mtv6w:
         (section==2'b10)? mtv7w:
                           mtv8w;
wire [79:0]         // error
  sumdata1w = sumdata1,                                                                                                                         
  sumdata2w = (layer_i==2'b00)? sumdata1:
              (layer_i==2'b01)? (rotat_en[1])?{sumdata1[59:0],sumdata1[79:60]} : {sumdata1[64:0],sumdata1[79:65]}:
              (layer_i==2'b10)? (rotat_en[1])?{sumdata1[9:0],sumdata1[79:10]} : {sumdata1[14:0],sumdata1[79:15]} :
                                (rotat_en[1])?{sumdata1[4:0],sumdata1[79:5]} : {sumdata1[9:0],sumdata1[79:10]}   ,
  sumdata3w = (layer_i==2'b00)? sumdata1:
              (layer_i==2'b01)? (rotat_en[2])?{sumdata1[19:0],sumdata1[79:20]} : {sumdata1[24:0],sumdata1[79:25]}:
              (layer_i==2'b10)? (rotat_en[2])?{sumdata1[39:0],sumdata1[79:40]} : {sumdata1[44:0],sumdata1[79:45]}:
                                (rotat_en[2])?{sumdata1[14:0],sumdata1[79:15]} : {sumdata1[19:0],sumdata1[79:20]},
  sumdata4w = (layer_i==2'b00)? sumdata1:
              (layer_i==2'b01)? (rotat_en[3])?{sumdata1[29:0],sumdata1[79:30]} : {sumdata1[34:0],sumdata1[79:35]}:
              (layer_i==2'b10)? (rotat_en[3])?{sumdata1[34:0],sumdata1[79:35]} : {sumdata1[39:0],sumdata1[79:40]}:
                                (rotat_en[3])?{sumdata1[9:0],sumdata1[79:10]} : {sumdata1[14:0],sumdata1[79:15]} ,
  sumdata5w = (layer_i==2'b00)? sumdata2:
              (layer_i==2'b01)? (rotat_en[4])?{sumdata2[69:0],sumdata2[79:70]} : {sumdata2[74:0],sumdata2[79:75]}:
              (layer_i==2'b10)? (rotat_en[4])?{sumdata2[44:0],sumdata2[79:45]} : {sumdata2[49:0],sumdata2[79:50]}:
                                (rotat_en[4])?{sumdata2[59:0],sumdata2[79:60]} : {sumdata2[64:0],sumdata2[79:65]},
  sumdata6w = (layer_i==2'b00)? sumdata2:
              (layer_i==2'b01)? (rotat_en[5])?{sumdata2[44:0],sumdata2[79:45]} : {sumdata2[49:0],sumdata2[79:50]}:
              (layer_i==2'b10)? (rotat_en[5])?{sumdata2[59:0],sumdata2[79:60]} : {sumdata2[64:0],sumdata2[79:65]}:
                                (rotat_en[5])? sumdata2  : {sumdata2[4:0],sumdata2[79:5]}                        ,
  sumdata7w = (layer_i==2'b00)? sumdata2:
              (layer_i==2'b01)? (rotat_en[6])?{sumdata2[14:0],sumdata2[79:15]} : {sumdata2[19:0],sumdata2[79:20]}:
              (layer_i==2'b10)? (rotat_en[6])?{sumdata2[9:0],sumdata2[79:10]} : {sumdata2[14:0],sumdata2[79:15]} :
                                (rotat_en[6])?{sumdata2[44:0],sumdata2[79:45]} : {sumdata2[49:0],sumdata2[79:50]},
  sumdata8w = (layer_i==2'b00)? sumdata2:
              (layer_i==2'b01)? (rotat_en[7])?{sumdata2[59:0],sumdata2[79:60]} : {sumdata2[64:0],sumdata2[79:65]}:
              (layer_i==2'b10)? (rotat_en[7])?{sumdata2[29:0],sumdata2[79:30]} : {sumdata2[34:0],sumdata2[79:35]}:
                                (rotat_en[7])? sumdata2 : {sumdata2[4:0],sumdata2[79:5]}                         ;

wire [79:0]
  sumdata1_w=(section==2'b00)? sumdata1w:
             (section==2'b01)? sumdata2w:
             (section==2'b10)? sumdata3w:
                               sumdata4w,
  sumdata2_w=(section==2'b00)? sumdata5w:
             (section==2'b01)? sumdata6w:
             (section==2'b10)? sumdata7w:
                               sumdata8w;
endmodule

module invpermutator2(
                      layer_i,section,
                      mtv1,mtv2,
                      mtv1_w,mtv2_w,
                      sumdata1,sumdata2,sumdata1_w,sumdata2_w,
                      rotat_en,
                      ctm1_i,ctm2_i,ctm1,ctm2);

input [1:0] layer_i,section;
input [79:0] mtv1,mtv2;
input [47:0] ctm1_i,ctm2_i;
input [79:0] sumdata1,sumdata2;
input [7:0]rotat_en;
output [47:0] ctm1,ctm2;
output [79:0] mtv1_w,mtv2_w;
output [79:0] sumdata1_w,sumdata2_w;
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//            2st row block   3st row block    4st row block
// shift Ext number  5             15           14
// shift Ext number  7             10           0
// shift Ext number  5             1            12
// shift Ext number  1             15           11
// shift Ext number  0             6            1
// shift Ext number  9             13           7
// shift Ext number  9             9            4
// shift Ext number  12            2            13
wire [47:0]
  ctm1_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[0])?{ctm1_i[17:0],ctm1_i[47:18]} : {ctm1_i[14:0],ctm1_i[47:15]} :
         (layer_i==2'b10)?(rotat_en[0])? ctm1_i : {ctm1_i[44:0],ctm1_i[47:45]} :
                          (rotat_en[0])?{ctm1_i[44:0],ctm1_i[47:45]} : {ctm1_i[41:0],ctm1_i[47:42]} ,
  ctm2_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[1])?{ctm1_i[23:0],ctm1_i[47:24]} : {ctm1_i[20:0],ctm1_i[47:21]} :
         (layer_i==2'b10)?(rotat_en[1])?{ctm1_i[32:0],ctm1_i[47:33]} : {ctm1_i[29:0],ctm1_i[47:30]} :
                          (rotat_en[1])?{ctm1_i[2:0],ctm1_i[47:3]} : ctm1_i ,
  ctm3_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[2])?{ctm1_i[17:0],ctm1_i[47:18]} : {ctm1_i[14:0],ctm1_i[47:15]} :
         (layer_i==2'b10)?(rotat_en[2])?{ctm1_i[5:0],ctm1_i[47:6]} : {ctm1_i[2:0],ctm1_i[47:3]} :
                          (rotat_en[2])?{ctm1_i[38:0],ctm1_i[47:39]} : {ctm1_i[35:0],ctm1_i[47:36]} ,
  ctm4_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[3])?{ctm1_i[5:0],ctm1_i[47:6]} : {ctm1_i[2:0],ctm1_i[47:3]} :
         (layer_i==2'b10)?(rotat_en[3])? ctm1_i : {ctm1_i[44:0],ctm1_i[47:45]} :
                          (rotat_en[3])?{ctm1_i[35:0],ctm1_i[47:36]} : {ctm1_i[32:0],ctm1_i[47:33]} ,
  ctm5_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[4])?{ctm2_i[2:0],ctm2_i[47:3]} : ctm2_i :
         (layer_i==2'b10)?(rotat_en[4])?{ctm2_i[20:0],ctm2_i[47:21]} : {ctm2_i[17:0],ctm2_i[47:18]} :
                          (rotat_en[4])?{ctm2_i[5:0],ctm2_i[47:6]} : {ctm2_i[2:0],ctm2_i[47:3]} ,
  ctm6_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[5])?{ctm2_i[29:0],ctm2_i[47:30]} : {ctm2_i[26:0],ctm2_i[47:27]} :
         (layer_i==2'b10)?(rotat_en[5])?{ctm2_i[41:0],ctm2_i[47:42]} : {ctm2_i[38:0],ctm2_i[47:39]} :
                          (rotat_en[5])?{ctm2_i[23:0],ctm2_i[47:24]} : {ctm2_i[20:0],ctm2_i[47:21]} ,
  ctm7_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[6])?{ctm2_i[29:0],ctm2_i[47:30]} : {ctm2_i[26:0],ctm2_i[47:27]} :
         (layer_i==2'b10)?(rotat_en[6])?{ctm2_i[29:0],ctm2_i[47:30]} : {ctm2_i[26:0],ctm2_i[47:27]} :
                          (rotat_en[6])?{ctm2_i[14:0],ctm2_i[47:15]} : {ctm2_i[11:0],ctm2_i[47:12]} ,
  ctm8_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[7])?{ctm2_i[38:0],ctm2_i[47:39]} : {ctm2_i[35:0],ctm2_i[47:36]} :
         (layer_i==2'b10)?(rotat_en[7])?{ctm2_i[8:0],ctm2_i[47:9]} : {ctm2_i[5:0],ctm2_i[47:6]} :
                          (rotat_en[7])?{ctm2_i[41:0],ctm2_i[47:42]} : {ctm2_i[38:0],ctm2_i[47:39]} ;
wire [47:0]
     ctm1=(section==2'b00)?ctm1_w:
          (section==2'b01)?ctm2_w:
          (section==2'b10)?ctm3_w:
                           ctm4_w,
     ctm2=(section==2'b00)?ctm5_w:
          (section==2'b01)?ctm6_w:
          (section==2'b10)?ctm7_w:
                           ctm8_w;

wire [79:0]
     mtv9w=  (layer_i==2'b00)? mtv1:
             (layer_i==2'b01)? (rotat_en[0])?{mtv1[49:0],mtv1[79:50]} : {mtv1[54:0],mtv1[79:55]}:
             (layer_i==2'b10)? (rotat_en[0])? mtv1: {mtv1[4:0],mtv1[79:5]}                       :
                               (rotat_en[0])?{mtv1[4:0],mtv1[79:5]} : {mtv1[9:0],mtv1[79:10]}   ,
     mtv10w= (layer_i==2'b00)? mtv1:
             (layer_i==2'b01)? (rotat_en[1])?{mtv1[39:0],mtv1[79:40]} : {mtv1[44:0],mtv1[79:45]}:
             (layer_i==2'b10)? (rotat_en[1])?{mtv1[24:0],mtv1[79:25]} : {mtv1[29:0],mtv1[79:30]}:
                               (rotat_en[1])?{mtv1[74:0],mtv1[79:75]} : mtv1,
     mtv11w= (layer_i==2'b00)? mtv1:
             (layer_i==2'b01)? (rotat_en[2])?{mtv1[49:0],mtv1[79:50]} : {mtv1[54:0],mtv1[79:55]}:
             (layer_i==2'b10)? (rotat_en[2])?{mtv1[69:0],mtv1[79:70]} : {mtv1[74:0],mtv1[79:75]}:
                               (rotat_en[2])?{mtv1[14:0],mtv1[79:15]} : {mtv1[19:0],mtv1[79:20]},
     mtv12w= (layer_i==2'b00)? mtv1:
             (layer_i==2'b01)? (rotat_en[3])?{mtv1[69:0],mtv1[79:70]} : {mtv1[74:0],mtv1[79:75]}:
             (layer_i==2'b10)? (rotat_en[3])? mtv1 : {mtv1[4:0],mtv1[79:5]}                      :
                               (rotat_en[3])?{mtv1[19:0],mtv1[79:20]} : {mtv1[24:0],mtv1[79:25]},
     mtv13w= (layer_i==2'b00)? mtv2:
             (layer_i==2'b01)? (rotat_en[4])?{mtv2[74:0],mtv2[79:75]}  : mtv2:
             (layer_i==2'b10)? (rotat_en[4])?{mtv2[44:0],mtv2[79:45]} : {mtv2[49:0],mtv2[79:50]}:
                               (rotat_en[4])?{mtv2[69:0],mtv2[79:70]} : {mtv2[74:0],mtv2[79:75]},
     mtv14w= (layer_i==2'b00)? mtv2:
             (layer_i==2'b01)? (rotat_en[5])?{mtv2[29:0],mtv2[79:30]} : {mtv2[34:0],mtv2[79:35]}:
             (layer_i==2'b10)? (rotat_en[5])?{mtv2[9:0],mtv2[79:10]} : {mtv2[14:0],mtv2[79:15]} :
                               (rotat_en[5])?{mtv2[39:0],mtv2[79:40]} : {mtv2[44:0],mtv2[79:45]},
     mtv15w= (layer_i==2'b00)? mtv2:
             (layer_i==2'b01)? (rotat_en[6])?{mtv2[29:0],mtv2[79:30]} : {mtv2[34:0],mtv2[79:35]}:
             (layer_i==2'b10)? (rotat_en[6])?{mtv2[29:0],mtv2[79:30]} : {mtv2[34:0],mtv2[79:35]}:
                               (rotat_en[6])?{mtv2[54:0],mtv2[79:55]} : {mtv2[59:0],mtv2[79:60]},
     mtv16w= (layer_i==2'b00)? mtv2:
             (layer_i==2'b01)? (rotat_en[7])?{mtv2[14:0],mtv2[79:15]} : {mtv2[19:0],mtv2[79:20]}:
             (layer_i==2'b10)? (rotat_en[7])?{mtv2[64:0],mtv2[79:65]} : {mtv2[69:0],mtv2[79:70]}:
                               (rotat_en[7])?{mtv2[9:0],mtv2[79:10]} : {mtv2[14:0],mtv2[79:15]} ;

wire [79:0]
  mtv1_w = (section==2'b00)? mtv9w:
           (section==2'b01)? mtv10w:
           (section==2'b10)? mtv11w:
                             mtv12w,
  mtv2_w= (section==2'b00)? mtv13w:
          (section==2'b01)? mtv14w:
          (section==2'b10)? mtv15w:
                            mtv16w;
wire [79:0]
     sumdata9w=  (layer_i==2'b00)? sumdata1:
                 (layer_i==2'b01)? (rotat_en[0])?{sumdata1[49:0],sumdata1[79:50]} : {sumdata1[54:0],sumdata1[79:55]}:
                 (layer_i==2'b10)? (rotat_en[0])? sumdata1: {sumdata1[4:0],sumdata1[79:5]}                          :
                                   (rotat_en[0])?{sumdata1[4:0],sumdata1[79:5]} : {sumdata1[9:0],sumdata1[79:10]}   ,
     sumdata10w= (layer_i==2'b00)? sumdata1:
                 (layer_i==2'b01)? (rotat_en[1])?{sumdata1[39:0],sumdata1[79:40]} : {sumdata1[44:0],sumdata1[79:45]}:
                 (layer_i==2'b10)? (rotat_en[1])?{sumdata1[24:0],sumdata1[79:25]} : {sumdata1[29:0],sumdata1[79:30]}:
                                   (rotat_en[1])?{sumdata1[74:0],sumdata1[79:75]} : sumdata1                          ,
     sumdata11w= (layer_i==2'b00)? sumdata1:
                 (layer_i==2'b01)? (rotat_en[2])?{sumdata1[49:0],sumdata1[79:50]} : {sumdata1[54:0],sumdata1[79:55]}:
                 (layer_i==2'b10)? (rotat_en[2])?{sumdata1[69:0],sumdata1[79:70]} : {sumdata1[74:0],sumdata1[79:75]}:
                                   (rotat_en[2])?{sumdata1[14:0],sumdata1[79:15]} : {sumdata1[19:0],sumdata1[79:20]},
     sumdata12w= (layer_i==2'b00)? sumdata1:
                 (layer_i==2'b01)? (rotat_en[3])?{sumdata1[69:0],sumdata1[79:70]} : {sumdata1[74:0],sumdata1[79:75]}:
                 (layer_i==2'b10)? (rotat_en[3])? sumdata1 : {sumdata1[4:0],sumdata1[79:5]}                         :
                                   (rotat_en[3])?{sumdata1[19:0],sumdata1[79:20]} : {sumdata1[24:0],sumdata1[79:25]},
     sumdata13w= (layer_i==2'b00)? sumdata2:
                 (layer_i==2'b01)? (rotat_en[4])?{sumdata2[74:0],sumdata2[79:75]}  : sumdata2                          :
                 (layer_i==2'b10)? (rotat_en[4])?{sumdata2[44:0],sumdata2[79:45]} : {sumdata2[49:0],sumdata2[79:50]}:
                                   (rotat_en[4])?{sumdata2[69:0],sumdata2[79:70]} : {sumdata2[74:0],sumdata2[79:75]},
     sumdata14w= (layer_i==2'b00)? sumdata2:
                 (layer_i==2'b01)? (rotat_en[5])?{sumdata2[29:0],sumdata2[79:30]} : {sumdata2[34:0],sumdata2[79:35]}:
                 (layer_i==2'b10)? (rotat_en[5])?{sumdata2[9:0],sumdata2[79:10]} : {sumdata2[14:0],sumdata2[79:15]} :
                                   (rotat_en[5])?{sumdata2[39:0],sumdata2[79:40]} : {sumdata2[44:0],sumdata2[79:45]},
     sumdata15w= (layer_i==2'b00)? sumdata2:
                 (layer_i==2'b01)? (rotat_en[6])?{sumdata2[29:0],sumdata2[79:30]} : {sumdata2[34:0],sumdata2[79:35]}:
                 (layer_i==2'b10)? (rotat_en[6])?{sumdata2[29:0],sumdata2[79:30]} : {sumdata2[34:0],sumdata2[79:35]}:
                                   (rotat_en[6])?{sumdata2[54:0],sumdata2[79:55]} : {sumdata2[59:0],sumdata2[79:60]},
     sumdata16w= (layer_i==2'b00)? sumdata2:
                 (layer_i==2'b01)? (rotat_en[7])?{sumdata2[14:0],sumdata2[79:15]} : {sumdata2[19:0],sumdata2[79:20]}:
                 (layer_i==2'b10)? (rotat_en[7])?{sumdata2[64:0],sumdata2[79:65]} : {sumdata2[69:0],sumdata2[79:70]}:
                                   (rotat_en[7])?{sumdata2[9:0],sumdata2[79:10]} : {sumdata2[14:0],sumdata2[79:15]} ;

wire [79:0]
  sumdata1_w = (section==2'b00)? sumdata9w:
               (section==2'b01)? sumdata10w:
               (section==2'b10)? sumdata11w:
                                 sumdata12w,
  sumdata2_w= (section==2'b00)? sumdata13w:
              (section==2'b01)? sumdata14w:
              (section==2'b10)? sumdata15w:
                                sumdata16w;
endmodule

module invpermutator3(
                   layer_i,section,
                   mtv1,mtv2,
                   mtv1_w,mtv2_w,
                   sumdata1,sumdata2,sumdata1_w,sumdata2_w,                                                                                     
                   rotat_en,
                   ctm1_i,ctm2_i,ctm1,ctm2);

input [1:0] layer_i,section;
input [79:0] mtv1,mtv2;
input [47:0] ctm1_i,ctm2_i;
input [79:0] sumdata1,sumdata2;
input [7:0]rotat_en;
output [47:0] ctm1,ctm2;
output [79:0] mtv1_w,mtv2_w;
output [79:0] sumdata1_w,sumdata2_w;
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//            2st row block   3st row block    4st row block
// shift Ext number 14               4             1
// shift Ext number 0                14            2
// shift Ext number 13               14            3
// shift Ext number 4                7             14
// shift Ext number 0                3             4
// shift Ext number 8                12            1
// shift Ext number 3                4             10
// shift Ext number 0                2             6
wire [47:0]
  ctm1_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[0])?{ctm1_i[44:0],ctm1_i[47:45]} : {ctm1_i[41:0],ctm1_i[47:42]} :
         (layer_i==2'b10)?(rotat_en[0])?{ctm1_i[14:0],ctm1_i[47:15]} : {ctm1_i[11:0],ctm1_i[47:12]} :
                          (rotat_en[0])?{ctm1_i[5:0],ctm1_i[47:6]} : {ctm1_i[2:0],ctm1_i[47:3]} ,
  ctm2_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[1])?{ctm1_i[2:0],ctm1_i[47:3]} : ctm1_i :
         (layer_i==2'b10)?(rotat_en[1])?{ctm1_i[44:0],ctm1_i[47:45]} : {ctm1_i[41:0],ctm1_i[47:42]} :
                          (rotat_en[1])?{ctm1_i[8:0],ctm1_i[47:9]} : {ctm1_i[5:0],ctm1_i[47:6]} ,
  ctm3_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[2])?{ctm1_i[41:0],ctm1_i[47:42]} : {ctm1_i[38:0],ctm1_i[47:39]} :
         (layer_i==2'b10)?(rotat_en[2])?{ctm1_i[44:0],ctm1_i[47:45]} : {ctm1_i[41:0],ctm1_i[47:42]} :
                          (rotat_en[2])?{ctm1_i[11:0],ctm1_i[47:12]} : {ctm1_i[8:0],ctm1_i[47:9]} ,
  ctm4_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[3])?{ctm1_i[14:0],ctm1_i[47:15]} : {ctm1_i[11:0],ctm1_i[47:12]} :
         (layer_i==2'b10)?(rotat_en[3])?{ctm1_i[23:0],ctm1_i[47:24]} : {ctm1_i[20:0],ctm1_i[47:21]} :
                          (rotat_en[3])?{ctm1_i[44:0],ctm1_i[47:45]} : {ctm1_i[41:0],ctm1_i[47:42]} ,
  ctm5_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?ctm2_i:
         (layer_i==2'b10)?(rotat_en[4])?{ctm2_i[11:0],ctm2_i[47:12]} : {ctm2_i[8:0],ctm2_i[47:9]} :
                          (rotat_en[4])?{ctm2_i[14:0],ctm2_i[47:15]} : {ctm2_i[11:0],ctm2_i[47:12]} ,
  ctm6_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[5])?{ctm2_i[26:0],ctm2_i[47:27]} : {ctm2_i[23:0],ctm2_i[47:24]} :
         (layer_i==2'b10)?(rotat_en[5])?{ctm2_i[38:0],ctm2_i[47:39]} : {ctm2_i[35:0],ctm2_i[47:36]} :
                          (rotat_en[5])?{ctm2_i[5:0],ctm2_i[47:6]} : {ctm2_i[2:0],ctm2_i[47:3]} ,
  ctm7_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[6])?{ctm2_i[11:0],ctm2_i[47:12]} : {ctm2_i[8:0],ctm2_i[47:9]} :
         (layer_i==2'b10)?(rotat_en[6])?{ctm2_i[14:0],ctm2_i[47:15]} : {ctm2_i[11:0],ctm2_i[47:12]} :
                          (rotat_en[6])?{ctm2_i[32:0],ctm2_i[47:33]} : {ctm2_i[29:0],ctm2_i[47:30]} ,
  ctm8_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[7])?{ctm2_i[2:0],ctm2_i[47:3]} : ctm2_i :
         (layer_i==2'b10)?(rotat_en[7])?{ctm2_i[8:0],ctm2_i[47:9]} : {ctm2_i[5:0],ctm2_i[47:6]} :
                          (rotat_en[7])?{ctm2_i[20:0],ctm2_i[47:21]} : {ctm2_i[17:0],ctm2_i[47:18]} ;
wire [47:0]
     ctm1=(section==2'b00)?ctm1_w:
          (section==2'b01)?ctm2_w:
          (section==2'b10)?ctm3_w:
                           ctm4_w,
     ctm2=(section==2'b00)?ctm5_w:
          (section==2'b01)?ctm6_w:
          (section==2'b10)?ctm7_w:
                           ctm8_w;
 //            2st row block   3st row block    4st row block
// shift Ext number 14               4             1
// shift Ext number 0                14            2
// shift Ext number 13               14            3
// shift Ext number 4                7             14
// shift Ext number 0                3             4
// shift Ext number 8                12            1
// shift Ext number 3                4             10
// shift Ext number 0                2             6
wire [79:0]
  mtv17w = (layer_i==2'b00)?  mtv1:
           (layer_i==2'b01)?  (rotat_en[0])?{mtv1[4:0],mtv1[79:5]} : {mtv1[9:0],mtv1[79:10]}   :
           (layer_i==2'b10)?  (rotat_en[0])?{mtv1[54:0],mtv1[79:55]} : {mtv1[59:0],mtv1[79:60]}:
                              (rotat_en[0])?{mtv1[69:0],mtv1[79:70]} : {mtv1[74:0],mtv1[79:75]},
  mtv18w = (layer_i==2'b00)?  mtv1:
           (layer_i==2'b01)?  (rotat_en[1])?{mtv1[74:0],mtv1[79:75]}  : mtv1                   :
           (layer_i==2'b10)?  (rotat_en[1])?{mtv1[4:0],mtv1[79:5]} : {mtv1[9:0],mtv1[79:10]}   :
                              (rotat_en[1])?{mtv1[64:0],mtv1[79:65]} : {mtv1[69:0],mtv1[79:70]},
  mtv19w = (layer_i==2'b00)?  mtv1:
           (layer_i==2'b01)?  (rotat_en[2])?{mtv1[9:0],mtv1[79:10]} : {mtv1[14:0],mtv1[79:15]} :
           (layer_i==2'b10)?  (rotat_en[2])?{mtv1[4:0],mtv1[79:5]} : {mtv1[9:0],mtv1[79:10]}   :
                              (rotat_en[2])?{mtv1[59:0],mtv1[79:60]} : {mtv1[64:0],mtv1[79:65]},
  mtv20w = (layer_i==2'b00)?  mtv1:
           (layer_i==2'b01)?  (rotat_en[3])?{mtv1[54:0],mtv1[79:55]} : {mtv1[59:0],mtv1[79:60]}:
           (layer_i==2'b10)?  (rotat_en[3])?{mtv1[39:0],mtv1[79:40]} : {mtv1[44:0],mtv1[79:45]}:
                              (rotat_en[3])?{mtv1[4:0],mtv1[79:5]} : {mtv1[9:0],mtv1[79:10]}   ,
  mtv21w = (layer_i==2'b00)?  mtv2:
           (layer_i==2'b01)?   mtv2:
           (layer_i==2'b10)?  (rotat_en[4])?{mtv2[59:0],mtv2[79:60]} : {mtv2[64:0],mtv2[79:65]}:
                              (rotat_en[4])?{mtv2[54:0],mtv2[79:55]} : {mtv2[59:0],mtv2[79:60]},
  mtv22w = (layer_i==2'b00)?  mtv2:
           (layer_i==2'b01)?  (rotat_en[5])?{mtv2[34:0],mtv2[79:35]} : {mtv2[39:0],mtv2[79:40]}:
           (layer_i==2'b10)?  (rotat_en[5])?{mtv2[14:0],mtv2[79:15]} : {mtv2[19:0],mtv2[79:20]}:
                              (rotat_en[5])?{mtv2[69:0],mtv2[79:70]} : {mtv2[74:0],mtv2[79:75]},
  mtv23w = (layer_i==2'b00)?  mtv2:
           (layer_i==2'b01)?  (rotat_en[6])?{mtv2[59:0],mtv2[79:60]} : {mtv2[64:0],mtv2[79:65]}:
           (layer_i==2'b10)?  (rotat_en[6])?{mtv2[54:0],mtv2[79:55]} : {mtv2[59:0],mtv2[79:60]}:
                              (rotat_en[6])?{mtv2[24:0],mtv2[79:25]} : {mtv2[29:0],mtv2[79:30]},
  mtv24w = (layer_i==2'b00)?  mtv2:
           (layer_i==2'b01)?  (rotat_en[7])?{mtv2[74:0],mtv2[79:75]}  : mtv2                   :
           (layer_i==2'b10)?  (rotat_en[7])?{mtv2[64:0],mtv2[79:65]} : {mtv2[69:0],mtv2[79:70]}:
                              (rotat_en[7])?{mtv2[44:0],mtv2[79:45]} : {mtv2[49:0],mtv2[79:50]};

wire [79:0]
  mtv1_w = (section==2'b00)? mtv17w :
           (section==2'b01)? mtv18w :
           (section==2'b10)? mtv19w :
                             mtv20w,
  mtv2_w = (section==2'b00)? mtv21w :
           (section==2'b01)? mtv22w :
           (section==2'b10)? mtv23w :
                             mtv24w;
wire [79:0]
  sumdata17w = (layer_i==2'b00)?  sumdata1:
               (layer_i==2'b01)?  (rotat_en[0])?{sumdata1[4:0],sumdata1[79:5]} : {sumdata1[9:0],sumdata1[79:10]}   :
               (layer_i==2'b10)?  (rotat_en[0])?{sumdata1[54:0],sumdata1[79:55]} : {sumdata1[59:0],sumdata1[79:60]}:
                                  (rotat_en[0])?{sumdata1[69:0],sumdata1[79:70]} : {sumdata1[74:0],sumdata1[79:75]},
  sumdata18w = (layer_i==2'b00)?  sumdata1:
               (layer_i==2'b01)?  (rotat_en[1])?{sumdata1[74:0],sumdata1[79:75]}  : sumdata1                          :
               (layer_i==2'b10)?  (rotat_en[1])?{sumdata1[4:0],sumdata1[79:5]} : {sumdata1[9:0],sumdata1[79:10]}   :
                                  (rotat_en[1])?{sumdata1[64:0],sumdata1[79:65]} : {sumdata1[69:0],sumdata1[79:70]},
  sumdata19w = (layer_i==2'b00)?  sumdata1:
               (layer_i==2'b01)?  (rotat_en[2])?{sumdata1[9:0],sumdata1[79:10]} : {sumdata1[14:0],sumdata1[79:15]} :
               (layer_i==2'b10)?  (rotat_en[2])?{sumdata1[4:0],sumdata1[79:5]} : {sumdata1[9:0],sumdata1[79:10]}   :
                                  (rotat_en[2])?{sumdata1[59:0],sumdata1[79:60]} : {sumdata1[64:0],sumdata1[79:65]},
  sumdata20w = (layer_i==2'b00)?  sumdata1:
               (layer_i==2'b01)?  (rotat_en[3])?{sumdata1[54:0],sumdata1[79:55]} : {sumdata1[59:0],sumdata1[79:60]}:
               (layer_i==2'b10)?  (rotat_en[3])?{sumdata1[39:0],sumdata1[79:40]} : {sumdata1[44:0],sumdata1[79:45]}:
                                  (rotat_en[3])?{sumdata1[4:0],sumdata1[79:5]} : {sumdata1[9:0],sumdata1[79:10]}   ,
  sumdata21w = (layer_i==2'b00)?  sumdata2:
               (layer_i==2'b01)?   sumdata2                                                               :
               (layer_i==2'b10)?  (rotat_en[4])?{sumdata2[59:0],sumdata2[79:60]} : {sumdata2[64:0],sumdata2[79:65]}:
                                  (rotat_en[4])?{sumdata2[54:0],sumdata2[79:55]} : {sumdata2[59:0],sumdata2[79:60]},
  sumdata22w = (layer_i==2'b00)?  sumdata2:
               (layer_i==2'b01)?  (rotat_en[5])?{sumdata2[34:0],sumdata2[79:35]} : {sumdata2[39:0],sumdata2[79:40]}:
               (layer_i==2'b10)?  (rotat_en[5])?{sumdata2[14:0],sumdata2[79:15]} : {sumdata2[19:0],sumdata2[79:20]}:
                                  (rotat_en[5])?{sumdata2[69:0],sumdata2[79:70]} : {sumdata2[74:0],sumdata2[79:75]},
  sumdata23w = (layer_i==2'b00)?  sumdata2:
               (layer_i==2'b01)?  (rotat_en[6])?{sumdata2[59:0],sumdata2[79:60]} : {sumdata2[64:0],sumdata2[79:65]}:
               (layer_i==2'b10)?  (rotat_en[6])?{sumdata2[54:0],sumdata2[79:55]} : {sumdata2[59:0],sumdata2[79:60]}:
                                  (rotat_en[6])?{sumdata2[24:0],sumdata2[79:25]} : {sumdata2[29:0],sumdata2[79:30]},
  sumdata24w = (layer_i==2'b00)?  sumdata2:
               (layer_i==2'b01)?  (rotat_en[7])?{sumdata2[74:0],sumdata2[79:75]}  : sumdata2                          :
               (layer_i==2'b10)?  (rotat_en[7])?{sumdata2[64:0],sumdata2[79:65]} : {sumdata2[69:0],sumdata2[79:70]}:
                                  (rotat_en[7])?{sumdata2[44:0],sumdata2[79:45]} : {sumdata2[49:0],sumdata2[79:50]};

wire [79:0]
  sumdata1_w = (section==2'b00)? sumdata17w :
               (section==2'b01)? sumdata18w :
               (section==2'b10)? sumdata19w :
                                 sumdata20w,
  sumdata2_w = (section==2'b00)? sumdata21w :
               (section==2'b01)? sumdata22w :
               (section==2'b10)? sumdata23w :
                                 sumdata24w;
endmodule

module invpermutator4(
                   layer_i,section,
                   mtv1,mtv2,
                   mtv1_w,mtv2_w,
                   sumdata1,sumdata2,sumdata1_w,sumdata2_w,                                                                                     
                   rotat_en,
                   ctm1_i,ctm2_i,ctm1,ctm2);

input [1:0] layer_i,section;
input [79:0] mtv1,mtv2;
input [47:0] ctm1_i,ctm2_i;
input [79:0] sumdata1,sumdata2;
input [7:0]rotat_en;
output [47:0] ctm1,ctm2;
output [79:0] mtv1_w,mtv2_w;
output [79:0] sumdata1_w,sumdata2_w;
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//            2st row block   3st row block    4st row block
// shift Ext number   0             8             3
// shift Ext number   13            4             2
// shift Ext number   13            7             3
// shift Ext number   12            8             0
// shift Ext number   6             4             2
// shift Ext number   2             15            2
// shift Ext number   11            9             14
// shift Ext number   13            10            7
wire [47:0]
  ctm1_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[0])?{ctm1_i[2:0],ctm1_i[47:3]} : ctm1_i :
         (layer_i==2'b10)?(rotat_en[0])?{ctm1_i[26:0],ctm1_i[47:27]} : {ctm1_i[23:0],ctm1_i[47:24]} :
                          (rotat_en[0])?{ctm1_i[11:0],ctm1_i[47:12]} : {ctm1_i[8:0],ctm1_i[47:9]} ,
  ctm2_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[1])?{ctm1_i[41:0],ctm1_i[47:42]} : {ctm1_i[38:0],ctm1_i[47:39]} :
         (layer_i==2'b10)?(rotat_en[1])?{ctm1_i[14:0],ctm1_i[47:15]} : {ctm1_i[11:0],ctm1_i[47:12]} :
                          (rotat_en[1])?{ctm1_i[8:0],ctm1_i[47:9]} : {ctm1_i[5:0],ctm1_i[47:6]} ,
  ctm3_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[2])?{ctm1_i[41:0],ctm1_i[47:42]} : {ctm1_i[38:0],ctm1_i[47:39]} :
         (layer_i==2'b10)?(rotat_en[2])?{ctm1_i[23:0],ctm1_i[47:24]} : {ctm1_i[20:0],ctm1_i[47:21]} :
                          (rotat_en[2])?{ctm1_i[11:0],ctm1_i[47:12]} : {ctm1_i[8:0],ctm1_i[47:9]} ,
  ctm4_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[3])?{ctm1_i[38:0],ctm1_i[47:39]} : {ctm1_i[35:0],ctm1_i[47:36]} :
         (layer_i==2'b10)?(rotat_en[3])?{ctm1_i[26:0],ctm1_i[47:27]} : {ctm1_i[23:0],ctm1_i[47:24]} :
                          (rotat_en[3])?{ctm1_i[2:0],ctm1_i[47:3]} : ctm1_i ,
  ctm5_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[4])?{ctm2_i[20:0],ctm2_i[47:21]} : {ctm2_i[17:0],ctm2_i[47:18]} :
         (layer_i==2'b10)?(rotat_en[4])?{ctm2_i[14:0],ctm2_i[47:15]} : {ctm2_i[11:0],ctm2_i[47:12]} :
                          (rotat_en[4])?{ctm2_i[8:0],ctm2_i[47:9]} : {ctm2_i[5:0],ctm2_i[47:6]} ,
  ctm6_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[5])?{ctm2_i[8:0],ctm2_i[47:9]} : {ctm2_i[5:0],ctm2_i[47:6]} :
         (layer_i==2'b10)?(rotat_en[5])? ctm2_i : {ctm2_i[44:0],ctm2_i[47:45]} :
                          (rotat_en[5])?{ctm2_i[8:0],ctm2_i[47:9]} : {ctm2_i[5:0],ctm2_i[47:6]} ,
  ctm7_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[6])?{ctm2_i[35:0],ctm2_i[47:36]} : {ctm2_i[32:0],ctm2_i[47:33]} :
         (layer_i==2'b10)?(rotat_en[6])?{ctm2_i[29:0],ctm2_i[47:30]} : {ctm2_i[26:0],ctm2_i[47:27]} :
                          (rotat_en[6])?{ctm2_i[44:0],ctm2_i[47:45]} : {ctm2_i[41:0],ctm2_i[47:42]} ,
  ctm8_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[7])?{ctm2_i[41:0],ctm2_i[47:42]} : {ctm2_i[38:0],ctm2_i[47:39]} :
         (layer_i==2'b10)?(rotat_en[7])?{ctm2_i[32:0],ctm2_i[47:33]} : {ctm2_i[29:0],ctm2_i[47:30]} :
                          (rotat_en[7])?{ctm2_i[23:0],ctm2_i[47:24]} : {ctm2_i[20:0],ctm2_i[47:21]} ;
wire [47:0]
     ctm1=(section==2'b00)?ctm1_w:
          (section==2'b01)?ctm2_w:
          (section==2'b10)?ctm3_w:
                           ctm4_w,
     ctm2=(section==2'b00)?ctm5_w:
          (section==2'b01)?ctm6_w:
          (section==2'b10)?ctm7_w:
                           ctm8_w;
//            2st row block   3st row block    4st row block
// shift Ext number   0             8             3
// shift Ext number   13            4             2
// shift Ext number   13            7             3
// shift Ext number   12            8             0
// shift Ext number   6             4             2
// shift Ext number   2             15            2
// shift Ext number   11            9             14
// shift Ext number   13            10            7
wire [79:0]
  mtv25w= (layer_i==2'b00)?  mtv1:
          (layer_i==2'b01)?  (rotat_en[0])?{mtv1[74:0],mtv1[79:75]}  : mtv1                :
          (layer_i==2'b10)?  (rotat_en[0])?{mtv1[34:0],mtv1[79:35]} : {mtv1[39:0],mtv1[79:40]}:
                             (rotat_en[0])?{mtv1[59:0],mtv1[79:60]} : {mtv1[64:0],mtv1[79:65]},
  mtv26w= (layer_i==2'b00)?  mtv1:
          (layer_i==2'b01)?  (rotat_en[1])?{mtv1[9:0],mtv1[79:10]} : {mtv1[14:0],mtv1[79:15]} :
          (layer_i==2'b10)?  (rotat_en[1])?{mtv1[54:0],mtv1[79:55]} : {mtv1[59:0],mtv1[79:60]}:
                             (rotat_en[1])?{mtv1[64:0],mtv1[79:65]} : {mtv1[69:0],mtv1[79:70]},
  mtv27w= (layer_i==2'b00)?  mtv1:
          (layer_i==2'b01)?  (rotat_en[2])?{mtv1[9:0],mtv1[79:10]} : {mtv1[14:0],mtv1[79:15]} :
          (layer_i==2'b10)?  (rotat_en[2])?{mtv1[39:0],mtv1[79:40]} : {mtv1[44:0],mtv1[79:45]}:
                             (rotat_en[2])?{mtv1[59:0],mtv1[79:60]} : {mtv1[64:0],mtv1[79:65]},
  mtv28w= (layer_i==2'b00)?  mtv1:
          (layer_i==2'b01)?  (rotat_en[3])?{mtv1[14:0],mtv1[79:15]} : {mtv1[19:0],mtv1[79:20]}:
          (layer_i==2'b10)?  (rotat_en[3])?{mtv1[34:0],mtv1[79:35]} : {mtv1[39:0],mtv1[79:40]}:
                             (rotat_en[3])?{mtv1[74:0],mtv1[79:75]}  : mtv1                   ,
  mtv29w= (layer_i==2'b00)?  mtv2:
          (layer_i==2'b01)?  (rotat_en[4])?{mtv2[44:0],mtv2[79:45]} : {mtv2[49:0],mtv2[79:50]}:
          (layer_i==2'b10)?  (rotat_en[4])?{mtv2[54:0],mtv2[79:55]} : {mtv2[59:0],mtv2[79:60]}:
                             (rotat_en[4])?{mtv2[64:0],mtv2[79:65]} : {mtv2[69:0],mtv2[79:70]},
  mtv30w= (layer_i==2'b00)?  mtv2:
          (layer_i==2'b01)?  (rotat_en[5])?{mtv2[64:0],mtv2[79:65]} : {mtv2[69:0],mtv2[79:70]}:
          (layer_i==2'b10)?  (rotat_en[5])? mtv2 : {mtv2[4:0],mtv2[79:5]}                     :
                             (rotat_en[5])?{mtv2[64:0],mtv2[79:65]} : {mtv2[69:0],mtv2[79:70]},
  mtv31w= (layer_i==2'b00)?  mtv2:
          (layer_i==2'b01)?  (rotat_en[6])?{mtv2[19:0],mtv2[79:20]} : {mtv2[24:0],mtv2[79:25]}:
          (layer_i==2'b10)?  (rotat_en[6])?{mtv2[29:0],mtv2[79:30]} : {mtv2[34:0],mtv2[79:35]}:
                             (rotat_en[6])?{mtv2[4:0],mtv2[79:5]} : {mtv2[9:0],mtv2[79:10]}   ,
  mtv32w= (layer_i==2'b00)?  mtv2:
          (layer_i==2'b01)?  (rotat_en[7])?{mtv2[9:0],mtv2[79:10]} : {mtv2[14:0],mtv2[79:15]} :
          (layer_i==2'b10)?  (rotat_en[7])?{mtv2[24:0],mtv2[79:25]} : {mtv2[29:0],mtv2[79:30]}:
                             (rotat_en[7])?{mtv2[39:0],mtv2[79:40]} : {mtv2[44:0],mtv2[79:45]};

wire [79:0]
  mtv1_w= (section==2'b00)? mtv25w:
          (section==2'b01)? mtv26w:
          (section==2'b10)? mtv27w:
                            mtv28w,
  mtv2_w= (section==2'b00)? mtv29w:
          (section==2'b01)? mtv30w:
          (section==2'b10)? mtv31w:
                            mtv32w;
wire [79:0]
  sumdata25w= (layer_i==2'b00)?  sumdata1:
              (layer_i==2'b01)?  (rotat_en[0])?{sumdata1[74:0],sumdata1[79:75]}  : sumdata1                :
              (layer_i==2'b10)?  (rotat_en[0])?{sumdata1[34:0],sumdata1[79:35]} : {sumdata1[39:0],sumdata1[79:40]}:
                                 (rotat_en[0])?{sumdata1[59:0],sumdata1[79:60]} : {sumdata1[64:0],sumdata1[79:65]},
  sumdata26w= (layer_i==2'b00)?  sumdata1:
              (layer_i==2'b01)?  (rotat_en[1])?{sumdata1[9:0],sumdata1[79:10]} : {sumdata1[14:0],sumdata1[79:15]} :
              (layer_i==2'b10)?  (rotat_en[1])?{sumdata1[54:0],sumdata1[79:55]} : {sumdata1[59:0],sumdata1[79:60]}:
                                 (rotat_en[1])?{sumdata1[64:0],sumdata1[79:65]} : {sumdata1[69:0],sumdata1[79:70]},
  sumdata27w= (layer_i==2'b00)?  sumdata1:
              (layer_i==2'b01)?  (rotat_en[2])?{sumdata1[9:0],sumdata1[79:10]} : {sumdata1[14:0],sumdata1[79:15]} :
              (layer_i==2'b10)?  (rotat_en[2])?{sumdata1[39:0],sumdata1[79:40]} : {sumdata1[44:0],sumdata1[79:45]}:
                                 (rotat_en[2])?{sumdata1[59:0],sumdata1[79:60]} : {sumdata1[64:0],sumdata1[79:65]},
  sumdata28w= (layer_i==2'b00)?  sumdata1:
              (layer_i==2'b01)?  (rotat_en[3])?{sumdata1[14:0],sumdata1[79:15]} : {sumdata1[19:0],sumdata1[79:20]}:
              (layer_i==2'b10)?  (rotat_en[3])?{sumdata1[34:0],sumdata1[79:35]} : {sumdata1[39:0],sumdata1[79:40]}:
                                 (rotat_en[3])?{sumdata1[74:0],sumdata1[79:75]}  : sumdata1                       ,
  sumdata29w= (layer_i==2'b00)?  sumdata2:
              (layer_i==2'b01)?  (rotat_en[4])?{sumdata2[44:0],sumdata2[79:45]} : {sumdata2[49:0],sumdata2[79:50]}:
              (layer_i==2'b10)?  (rotat_en[4])?{sumdata2[54:0],sumdata2[79:55]} : {sumdata2[59:0],sumdata2[79:60]}:
                                 (rotat_en[4])?{sumdata2[64:0],sumdata2[79:65]} : {sumdata2[69:0],sumdata2[79:70]},
  sumdata30w= (layer_i==2'b00)?  sumdata2:
              (layer_i==2'b01)?  (rotat_en[5])?{sumdata2[64:0],sumdata2[79:65]} : {sumdata2[69:0],sumdata2[79:70]}:
              (layer_i==2'b10)?  (rotat_en[5])? sumdata2 : {sumdata2[4:0],sumdata2[79:5]}                         :
                                 (rotat_en[5])?{sumdata2[64:0],sumdata2[79:65]} : {sumdata2[69:0],sumdata2[79:70]},
  sumdata31w= (layer_i==2'b00)?  sumdata2:
              (layer_i==2'b01)?  (rotat_en[6])?{sumdata2[19:0],sumdata2[79:20]} : {sumdata2[24:0],sumdata2[79:25]}:
              (layer_i==2'b10)?  (rotat_en[6])?{sumdata2[29:0],sumdata2[79:30]} : {sumdata2[34:0],sumdata2[79:35]}:
                                 (rotat_en[6])?{sumdata2[4:0],sumdata2[79:5]} : {sumdata2[9:0],sumdata2[79:10]}   ,
  sumdata32w= (layer_i==2'b00)?  sumdata2:
              (layer_i==2'b01)?  (rotat_en[7])?{sumdata2[9:0],sumdata2[79:10]} : {sumdata2[14:0],sumdata2[79:15]} :
              (layer_i==2'b10)?  (rotat_en[7])?{sumdata2[24:0],sumdata2[79:25]} : {sumdata2[29:0],sumdata2[79:30]}:
                                 (rotat_en[7])?{sumdata2[39:0],sumdata2[79:40]} : {sumdata2[44:0],sumdata2[79:45]};

wire [79:0]
  sumdata1_w= (section==2'b00)? sumdata25w:
              (section==2'b01)? sumdata26w:
              (section==2'b10)? sumdata27w:
                                sumdata28w,
  sumdata2_w= (section==2'b00)? sumdata29w:
              (section==2'b01)? sumdata30w:
              (section==2'b10)? sumdata31w:
                                sumdata32w;
endmodule

module invpermutator5(
                   layer_i,section,
                   mtv1,mtv2,
                   mtv1_w,mtv2_w,
                   sumdata1,sumdata2,sumdata1_w,sumdata2_w,                                                                                     
                   rotat_en,
                   ctm1_i,ctm2_i,ctm1,ctm2);

input [1:0] layer_i;
input [1:0] section;
input [79:0] mtv1,mtv2;
input [47:0] ctm1_i,ctm2_i;
input [79:0] sumdata1,sumdata2;
input [7:0]rotat_en;
output [47:0] ctm1,ctm2;
output [79:0] mtv1_w,mtv2_w;
output [79:0] sumdata1_w,sumdata2_w;
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//  1st row block circulant=0
//            2st row block   3st row block    4st row block
// shift Ext number  11          11              11
// shift Ext number  4           13              14
// shift Ext number  10          0               12
// shift Ext number  5           5               6
// shift Ext number  3           2               12
// shift Ext number  3           0               7
// shift Ext number  4           1               8
// shift Ext number  8           10              6
wire [47:0]
  ctm1_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[0])?{ctm1_i[35:0],ctm1_i[47:36]} : {ctm1_i[32:0],ctm1_i[47:33]} :
         (layer_i==2'b10)?(rotat_en[0])?{ctm1_i[35:0],ctm1_i[47:36]} : {ctm1_i[32:0],ctm1_i[47:33]} :
                          (rotat_en[0])?{ctm1_i[35:0],ctm1_i[47:36]} : {ctm1_i[32:0],ctm1_i[47:33]} ,
  ctm2_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[1])?{ctm1_i[14:0],ctm1_i[47:15]} : {ctm1_i[11:0],ctm1_i[47:12]} :
         (layer_i==2'b10)?(rotat_en[1])?{ctm1_i[41:0],ctm1_i[47:42]} : {ctm1_i[38:0],ctm1_i[47:39]} :
                          (rotat_en[1])?{ctm1_i[44:0],ctm1_i[47:45]} : {ctm1_i[41:0],ctm1_i[47:42]} ,
  ctm3_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[2])?{ctm1_i[32:0],ctm1_i[47:33]} : {ctm1_i[29:0],ctm1_i[47:30]} :
         (layer_i==2'b10)?(rotat_en[2])?{ctm1_i[2:0],ctm1_i[47:3]} : ctm1_i :
                          (rotat_en[2])?{ctm1_i[38:0],ctm1_i[47:39]} : {ctm1_i[35:0],ctm1_i[47:36]} ,
  ctm4_w=(layer_i==2'b00)?ctm1_i:
         (layer_i==2'b01)?(rotat_en[3])?{ctm1_i[17:0],ctm1_i[47:18]} : {ctm1_i[14:0],ctm1_i[47:15]} :
         (layer_i==2'b10)?(rotat_en[3])?{ctm1_i[17:0],ctm1_i[47:18]} : {ctm1_i[14:0],ctm1_i[47:15]} :
                          (rotat_en[3])?{ctm1_i[20:0],ctm1_i[47:21]} : {ctm1_i[17:0],ctm1_i[47:18]} ,
  ctm5_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[4])?{ctm2_i[11:0],ctm2_i[47:12]} : {ctm2_i[8:0],ctm2_i[47:9]} :
         (layer_i==2'b10)?(rotat_en[4])?{ctm2_i[8:0],ctm2_i[47:9]} : {ctm2_i[5:0],ctm2_i[47:6]} :
                          (rotat_en[4])?{ctm2_i[38:0],ctm2_i[47:39]} : {ctm2_i[35:0],ctm2_i[47:36]} ,
  ctm6_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[5])?{ctm2_i[11:0],ctm2_i[47:12]} : {ctm2_i[8:0],ctm2_i[47:9]} :
         (layer_i==2'b10)?(rotat_en[5])?{ctm2_i[2:0],ctm2_i[47:3]} : ctm2_i :
                          (rotat_en[5])?{ctm2_i[23:0],ctm2_i[47:24]} : {ctm2_i[20:0],ctm2_i[47:21]} ,
  ctm7_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[6])?{ctm2_i[14:0],ctm2_i[47:15]} : {ctm2_i[11:0],ctm2_i[47:12]} :
         (layer_i==2'b10)?(rotat_en[6])?{ctm2_i[5:0],ctm2_i[47:6]} : {ctm2_i[2:0],ctm2_i[47:3]} :
                          (rotat_en[6])?{ctm2_i[26:0],ctm2_i[47:27]} : {ctm2_i[23:0],ctm2_i[47:24]} ,
  ctm8_w=(layer_i==2'b00)?ctm2_i:
         (layer_i==2'b01)?(rotat_en[7])?{ctm2_i[26:0],ctm2_i[47:27]} : {ctm2_i[23:0],ctm2_i[47:24]} :
         (layer_i==2'b10)?(rotat_en[7])?{ctm2_i[32:0],ctm2_i[47:33]} : {ctm2_i[29:0],ctm2_i[47:30]} :
                          (rotat_en[7])?{ctm2_i[20:0],ctm2_i[47:21]} : {ctm2_i[17:0],ctm2_i[47:18]} ;
wire [47:0]
     ctm1=(section==2'b00)?ctm1_w:
          (section==2'b01)?ctm2_w:
          (section==2'b10)?ctm3_w:
                           ctm4_w,
     ctm2=(section==2'b00)?ctm5_w:
          (section==2'b01)?ctm6_w:
          (section==2'b10)?ctm7_w:
                           ctm8_w;
//            2st row block   3st row block    4st row block
// shift Ext number    11          11              11
// shift Ext number    4           13              14
// shift Ext number    10          0               12
// shift Ext number    5           5               6
// shift Ext number    3           2               12
// shift Ext number    3           0               7
// shift Ext number    4           1               8
// shift Ext number    8           10              6
wire [79:0]
  mtv33w= (layer_i==2'b00)? mtv1:
          (layer_i==2'b01)? (rotat_en[0])?{mtv1[19:0],mtv1[79:20]} : {mtv1[24:0],mtv1[79:25]}:
          (layer_i==2'b10)? (rotat_en[0])?{mtv1[19:0],mtv1[79:20]} : {mtv1[24:0],mtv1[79:25]}:
                            (rotat_en[0])?{mtv1[19:0],mtv1[79:20]} : {mtv1[24:0],mtv1[79:25]},
  mtv34w= (layer_i==2'b00)? mtv1:
          (layer_i==2'b01)? (rotat_en[1])?{mtv1[54:0],mtv1[79:55]} : {mtv1[59:0],mtv1[79:60]}:
          (layer_i==2'b10)? (rotat_en[1])?{mtv1[9:0],mtv1[79:10]} : {mtv1[14:0],mtv1[79:15]} :
                            (rotat_en[1])?{mtv1[4:0],mtv1[79:5]} : {mtv1[9:0],mtv1[79:10]}   ,
  mtv35w= (layer_i==2'b00)? mtv1:
          (layer_i==2'b01)? (rotat_en[2])?{mtv1[24:0],mtv1[79:25]} : {mtv1[29:0],mtv1[79:30]}:
          (layer_i==2'b10)? (rotat_en[2])?{mtv1[74:0],mtv1[79:75]}  : mtv1                   :
                            (rotat_en[2])?{mtv1[14:0],mtv1[79:15]} : {mtv1[19:0],mtv1[79:20]},
  mtv36w= (layer_i==2'b00)? mtv1:
          (layer_i==2'b01)? (rotat_en[3])?{mtv1[49:0],mtv1[79:50]} : {mtv1[54:0],mtv1[79:55]}:
          (layer_i==2'b10)? (rotat_en[3])?{mtv1[49:0],mtv1[79:50]} : {mtv1[54:0],mtv1[79:55]}:
                            (rotat_en[3])?{mtv1[44:0],mtv1[79:45]} : {mtv1[49:0],mtv1[79:50]},
  mtv37w= (layer_i==2'b00)? mtv2:
          (layer_i==2'b01)? (rotat_en[4])?{mtv2[59:0],mtv2[79:60]} : {mtv2[64:0],mtv2[79:65]}:
          (layer_i==2'b10)? (rotat_en[4])?{mtv2[64:0],mtv2[79:65]} : {mtv2[69:0],mtv2[79:70]}:
                            (rotat_en[4])?{mtv2[14:0],mtv2[79:15]} : {mtv2[19:0],mtv2[79:20]},
  mtv38w= (layer_i==2'b00)? mtv2:
          (layer_i==2'b01)? (rotat_en[5])?{mtv2[59:0],mtv2[79:60]} : {mtv2[64:0],mtv2[79:65]}:
          (layer_i==2'b10)? (rotat_en[5])?{mtv2[74:0],mtv2[79:75]} : mtv2                    :
                            (rotat_en[5])?{mtv2[39:0],mtv2[79:40]} : {mtv2[44:0],mtv2[79:45]},
  mtv39w= (layer_i==2'b00)? mtv2:
          (layer_i==2'b01)? (rotat_en[6])?{mtv2[54:0],mtv2[79:55]} : {mtv2[59:0],mtv2[79:60]}:
          (layer_i==2'b10)? (rotat_en[6])?{mtv2[69:0],mtv2[79:70]} : {mtv2[74:0],mtv2[79:75]}:
                            (rotat_en[6])?{mtv2[34:0],mtv2[79:35]} : {mtv2[39:0],mtv2[79:40]},
  mtv40w= (layer_i==2'b00)? mtv2:
          (layer_i==2'b01)? (rotat_en[7])?{mtv2[34:0],mtv2[79:35]} : {mtv2[39:0],mtv2[79:40]}:
          (layer_i==2'b10)? (rotat_en[7])?{mtv2[24:0],mtv2[79:25]} : {mtv2[29:0],mtv2[79:30]}:
                            (rotat_en[7])?{mtv2[44:0],mtv2[79:45]} : {mtv2[49:0],mtv2[79:50]};

wire [79:0]
  mtv1_w= (section==2'b00)? mtv33w:
          (section==2'b01)? mtv34w:
          (section==2'b10)? mtv35w:
                            mtv36w,
  mtv2_w= (section==2'b00)? mtv37w:
          (section==2'b01)? mtv38w:
          (section==2'b10)? mtv39w:
                            mtv40w;
wire [79:0]
  sumdata33w= (layer_i==2'b00)? sumdata1:                                                                                                       
              (layer_i==2'b01)? (rotat_en[0])?{sumdata1[19:0],sumdata1[79:20]} : {sumdata1[24:0],sumdata1[79:25]}:
              (layer_i==2'b10)? (rotat_en[0])?{sumdata1[19:0],sumdata1[79:20]} : {sumdata1[24:0],sumdata1[79:25]}:
                                (rotat_en[0])?{sumdata1[19:0],sumdata1[79:20]} : {sumdata1[24:0],sumdata1[79:25]},
  sumdata34w= (layer_i==2'b00)? sumdata1:
              (layer_i==2'b01)? (rotat_en[1])?{sumdata1[54:0],sumdata1[79:55]} : {sumdata1[59:0],sumdata1[79:60]}:
              (layer_i==2'b10)? (rotat_en[1])?{sumdata1[9:0],sumdata1[79:10]} : {sumdata1[14:0],sumdata1[79:15]} :
                                (rotat_en[1])?{sumdata1[4:0],sumdata1[79:5]} : {sumdata1[9:0],sumdata1[79:10]}   ,
  sumdata35w= (layer_i==2'b00)? sumdata1:
              (layer_i==2'b01)? (rotat_en[2])?{sumdata1[24:0],sumdata1[79:25]} : {sumdata1[29:0],sumdata1[79:30]}:
              (layer_i==2'b10)? (rotat_en[2])?{sumdata1[74:0],sumdata1[79:75]}  : sumdata1                          :
                                (rotat_en[2])?{sumdata1[14:0],sumdata1[79:15]} : {sumdata1[19:0],sumdata1[79:20]},
  sumdata36w= (layer_i==2'b00)? sumdata1:
              (layer_i==2'b01)? (rotat_en[3])?{sumdata1[49:0],sumdata1[79:50]} : {sumdata1[54:0],sumdata1[79:55]}:
              (layer_i==2'b10)? (rotat_en[3])?{sumdata1[49:0],sumdata1[79:50]} : {sumdata1[54:0],sumdata1[79:55]}:
                                (rotat_en[3])?{sumdata1[44:0],sumdata1[79:45]} : {sumdata1[49:0],sumdata1[79:50]},
  sumdata37w= (layer_i==2'b00)? sumdata2:
              (layer_i==2'b01)? (rotat_en[4])?{sumdata2[59:0],sumdata2[79:60]} : {sumdata2[64:0],sumdata2[79:65]}:
              (layer_i==2'b10)? (rotat_en[4])?{sumdata2[64:0],sumdata2[79:65]} : {sumdata2[69:0],sumdata2[79:70]}:
                                (rotat_en[4])?{sumdata2[14:0],sumdata2[79:15]} : {sumdata2[19:0],sumdata2[79:20]},
  sumdata38w= (layer_i==2'b00)? sumdata2:
              (layer_i==2'b01)? (rotat_en[5])?{sumdata2[59:0],sumdata2[79:60]} : {sumdata2[64:0],sumdata2[79:65]}:
              (layer_i==2'b10)? (rotat_en[5])?{sumdata2[74:0],sumdata2[79:75]} : sumdata2                          :
                                (rotat_en[5])?{sumdata2[39:0],sumdata2[79:40]} : {sumdata2[44:0],sumdata2[79:45]},
  sumdata39w= (layer_i==2'b00)? sumdata2:
              (layer_i==2'b01)? (rotat_en[6])?{sumdata2[54:0],sumdata2[79:55]} : {sumdata2[59:0],sumdata2[79:60]}:
              (layer_i==2'b10)? (rotat_en[6])?{sumdata2[69:0],sumdata2[79:70]} : {sumdata2[74:0],sumdata2[79:75]}:
                                (rotat_en[6])?{sumdata2[34:0],sumdata2[79:35]} : {sumdata2[39:0],sumdata2[79:40]},
  sumdata40w= (layer_i==2'b00)? sumdata2:
              (layer_i==2'b01)? (rotat_en[7])?{sumdata2[34:0],sumdata2[79:35]} : {sumdata2[39:0],sumdata2[79:40]}:
              (layer_i==2'b10)? (rotat_en[7])?{sumdata2[24:0],sumdata2[79:25]} : {sumdata2[29:0],sumdata2[79:30]}:
                                (rotat_en[7])?{sumdata2[44:0],sumdata2[79:45]} : {sumdata2[49:0],sumdata2[79:50]};

wire [79:0]
  sumdata1_w= (section==2'b00)? sumdata33w:
              (section==2'b01)? sumdata34w:
              (section==2'b10)? sumdata35w:
                                sumdata36w,
  sumdata2_w= (section==2'b00)? sumdata37w:
              (section==2'b01)? sumdata38w:
              (section==2'b10)? sumdata39w:
                                sumdata40w;
endmodule

module controller(
                 RESET_N,CLK,
                 tmn,start_ldpc,start_Ldata,maxiter,
                 data_wrsa,data_wrsb,deca_en,decb_en,hb_en,load_data_en,
                 vncn_en,memwra_en,memwrb_en,dec_fin,hb_vlid,hboutmux,
                 layer_i,section,section_r,
                 iter_count,
                 vncn_count,
                 ch_counta,ch_countb,
                 addr_count,addr_ch_count,
                 hb_count,hb_count_wr,
                 memgroup_hb,section_hb);

input        RESET_N,CLK;
input        tmn,start_ldpc,start_Ldata;
input [4:0]  maxiter;
output       data_wrsa,data_wrsb,deca_en,decb_en,hb_en,load_data_en,
             vncn_en,memwra_en,memwrb_en,dec_fin,hb_vlid,hboutmux;
output [1:0]  layer_i,section,section_r;
output [4:0]  iter_count;
output [3:0]  vncn_count;
output [12:0] ch_counta,ch_countb;
output [3:0]  addr_count,addr_ch_count;
output [3:0]  hb_count,hb_count_wr;
output [2:0] memgroup_hb;
output [1:0] section_hb;
reg        data_wrsa,data_wrsb,hb_en,load_data_en,
           memwra_en,memwrb_en,dec_fin,hb_vlid;
reg [2:0]  state;
reg [3:0]  vncn_count;
reg [3:0]  addr_count,addr_ch_count;
reg [3:0]  hb_count,hb_count_wr;
reg [12:0] ch_counta,ch_countb;
reg [1:0]  layer_i,section,section_r;
reg [4:0]  iter_count;
reg [5:0]  memid_hb;
reg [2:0]  memgroup_hb;
reg [1:0]  section_hb;
parameter idle=3'b000,load_data=3'b001,
          dec_LdataB=3'b011,dec_LdataA=3'b100,hb_dec_LdataB=3'b101,
          hb_act=3'b111;
wire vncn_en=(state==dec_LdataB |
              state==dec_LdataA |
              state==hb_dec_LdataB ) & (vncn_count==4'd0);
wire deca_en=(state==dec_LdataB |
              state==hb_dec_LdataB) & (~(iter_count==maxiter));
wire decb_en=(state==dec_LdataA) & (~(iter_count==maxiter));
wire        hboutmux=(memid_hb==6'd1  | memid_hb==6'd3  | memid_hb==6'd5  |
                      memid_hb==6'd7  | memid_hb==6'd9   );
always @(negedge RESET_N or posedge CLK)
begin
  if (~RESET_N)
  begin
    state       <=0;
    data_wrsa   <=0;
    data_wrsb   <=0;
    hb_en       <=0;
    load_data_en<=0;
    memwra_en   <=0;
    memwrb_en   <=0;
    vncn_count  <=0;
    addr_count  <=0;
    addr_ch_count<=0;
    ch_counta   <=0;
    ch_countb   <=0;
    hb_count    <=0;
    layer_i     <=0;
    section     <=0;
    iter_count  <=0;
    dec_fin     <=1;
    hb_vlid     <=0;
    hb_count_wr <=0;
    memid_hb    <=0;
    memgroup_hb <=0;
    section_hb  <=0;
    section_r   <=0;
  end
  else
  begin
  section_r<=section;
    case(state)
      idle:
      begin
        hb_en       <=0;
        load_data_en<=0;
        memwra_en   <=0;
        memwrb_en   <=0;
        vncn_count  <=0;
        addr_count  <=0;
        addr_ch_count<=0;
        ch_counta   <=0;
        ch_countb   <=0;
        hb_count    <=0;
        layer_i     <=0;
        section     <=0;
        iter_count  <=0;
        data_wrsa   <=start_ldpc;
        data_wrsb   <=0;
        state       <=(start_ldpc)?load_data:idle;
        dec_fin     <=1;
        hb_vlid     <=0;
        hb_count_wr <=0;
        memid_hb    <=0;
        memgroup_hb <=0;
        section_hb  <=0;
      end
      load_data:
      begin
        data_wrsa   <=(ch_counta <13'd655);
        data_wrsb   <=0;
        hb_en       <=0;
        ch_counta   <=(ch_counta==13'd655)?13'd655:ch_counta+13'd1;
        ch_countb   <=0;
        hb_count    <=0;
        iter_count  <=0;
        load_data_en<=(ch_counta >=13'd15 );
        memwra_en   <=(ch_counta <13'd655);
        state       <=(ch_counta==13'd655)?dec_LdataB:load_data;
        memwrb_en   <=0;
        vncn_count  <=0;
        addr_count  <=0;
        addr_ch_count<=(addr_ch_count==4'd15 | ~data_wrsa)?4'd0:addr_ch_count+4'd1;
        layer_i     <=0;
        section     <=0;
        dec_fin     <=1;
        hb_vlid     <=0;
        hb_count_wr <=0;
        memid_hb    <=0;
        memgroup_hb <=0;
        section_hb  <=0;
      end
      dec_LdataB://state:4'b0011
      begin
        data_wrsa    <=(ch_countb==maxiter*768);
        data_wrsb    <=(ch_countb < 13'd656);
        load_data_en <=(ch_countb > 13'd15 & ch_countb < 13'd656);
        ch_counta    <=0;
        ch_countb    <=(ch_countb==maxiter*768)?13'd0:ch_countb+13'd1;
        addr_ch_count<=(ch_countb==13'd656 | addr_ch_count==4'd15 | ~data_wrsb)?4'd0:addr_ch_count+4'd1;
        hb_vlid      <=0;
        hb_en        <=0;
        hb_count     <=(hb_en)?(hb_count==4'd15)?4'd0:hb_count+4'd1:4'd0;
        memid_hb     <=0;
        memgroup_hb  <=0;
        section_hb   <=0;
        if(ch_countb==maxiter*768)
        begin
          state      <=(start_ldpc)?dec_LdataA:hb_act;
          memwra_en  <=0;
          memwrb_en  <=0;
          vncn_count <=0;
          addr_count <=0;
          layer_i    <=0;
          section    <=0;
          iter_count <=0;
          dec_fin    <=1;
          hb_count_wr<=0;
        end
        else
        begin
          state       <=dec_LdataB;
          memwra_en   <=(vncn_count==4'd4 | vncn_count==4'd6 | vncn_count==4'd8 | vncn_count==4'd10) ;
          memwrb_en   <=(ch_countb < 13'd656);
          if(layer_i==2'd3 & addr_count==4'd15 & vncn_count==4'd11 & section==2'd3)
            iter_count<=(iter_count==maxiter)?5'd8:iter_count +5'd1;
          if(addr_count==4'd15 & section==2'd3 & vncn_count==4'd11)
            layer_i   <=layer_i+2'd1;
          section     <=(vncn_count>=4'd4)? (~memwra_en)? section:section+2'd1:section+2'd1;
          addr_count  <=(section==2'd3 & vncn_count==4'd11)?addr_count+4'd1:addr_count;
          vncn_count  <=(vncn_count==4'd11)?4'd0:vncn_count+4'd1;
          dec_fin     <=0;
          hb_count_wr <=(section==2'd3 & vncn_count==4'd11)?hb_count_wr+4'd1:hb_count_wr;
        end
      end
      dec_LdataA://load sa data and hb sa output  state:4'b0100
      begin
        data_wrsa   <=(ch_counta <13'd656);
        data_wrsb   <=(ch_counta==maxiter*768-1);
        load_data_en<=(ch_counta >= 13'd15 & ch_counta < 13'd655);
        ch_counta   <=(ch_counta==maxiter*768-1)?13'd0:ch_counta+13'd1;
        ch_countb   <=0;
        hb_vlid     <=(ch_counta >=13'd17 & ch_counta <13'd657);
        hb_en       <=(ch_counta <13'd657);
        addr_ch_count<=(ch_counta==13'd656 | addr_ch_count==4'd15 | ~data_wrsa)?4'd0:addr_ch_count+4'd1;
        if(ch_counta==maxiter*768-1)
        begin
          state     <=(start_ldpc)?hb_dec_LdataB:hb_act;
          memwra_en <=0;
          memwrb_en <=0;
          vncn_count<=0;
          addr_count<=0;
          layer_i   <=0;
          section   <=0;
          iter_count<=0;
          hb_count  <=0;
          dec_fin   <=1;
          hb_count_wr <=0;
          memid_hb     <=0;
          memgroup_hb  <=0;
          section_hb   <=0;
        end
        else
        begin
          state       <=dec_LdataA;
          memwra_en   <=(ch_counta < 13'd656);
          memwrb_en   <=(vncn_count==4'd4 | vncn_count==4'd6 | vncn_count==4'd8 | vncn_count==4'd10) ;
          if(layer_i==2'd3 & addr_count==4'd15 & vncn_count==4'd11 & section==2'd3)
            iter_count<=(iter_count==maxiter)?5'd8:iter_count +5'd1;
          if(addr_count==4'd15 & section==2'd3 & vncn_count==4'd11)
            layer_i   <=layer_i+2'd1;
          section     <=(vncn_count>=4'd4)? (~memwrb_en)? section:section+2'd1:section+2'd1;
          addr_count  <=(section==2'd3 & vncn_count==4'd11)?addr_count+4'd1:addr_count;
          vncn_count  <=(vncn_count==4'd11)?4'd0:vncn_count+4'd1;
          hb_count    <=(hb_en)?(hb_count==4'd15)?4'd0:hb_count+4'd1:4'd0;
          dec_fin     <=0;
          hb_count_wr <=(section==2'd3 & vncn_count==4'd11)?hb_count_wr+4'd1:hb_count_wr;
          section_hb<=(hb_en)?((hb_count==4'd15)?
                       section_hb+2'd1:section_hb):2'd0 ;
          if(hb_vlid)
          begin
            if((hb_count==4'd0) & section_hb==2'd0)
              memid_hb<=(memid_hb==6'd15)? 6'd0 :
                     (~data_wrsa & ~data_wrsb)? 6'd0 : memid_hb+6'd1;
            if((memid_hb==6'd1 | memid_hb==6'd3 | memid_hb==6'd5 | memid_hb==6'd7 | memid_hb==6'd9) & (hb_count==4'd0) & section_hb==2'd0)
              memgroup_hb<=(memgroup_hb==3'd4)?
                         3'd0 : memgroup_hb+3'd1;
          end
        end
      end
      hb_dec_LdataB://state:4'b0101
      begin
        data_wrsa   <=(ch_countb==maxiter*768-1);
        data_wrsb   <=(ch_countb <13'd656);
        load_data_en<=(ch_countb>=13'd15 & ch_countb < 13'd655);
        ch_counta   <=0;
        ch_countb   <=(ch_countb==maxiter*768-1)?13'd0:ch_countb+13'd1;
        addr_ch_count<=(ch_countb==13'd656 | addr_ch_count==4'd15 | ~data_wrsb)?4'd0:addr_ch_count+4'd1;
        hb_vlid      <=(ch_countb >=13'd17 & ch_countb <13'd657);
        hb_en        <=(ch_countb <13'd656);
        if(ch_countb==maxiter*768-1)
        begin
          state     <=(start_ldpc)?dec_LdataA:hb_act;
          memwra_en <=0;
          memwrb_en <=0;
          vncn_count<=0;
          addr_count<=0;
          layer_i   <=0;
          section   <=0;
          iter_count<=0;
          hb_count  <=0;
          dec_fin   <=1;
          hb_count_wr<=0;
          memid_hb   <=0;
          memgroup_hb<=0;
          section_hb <=0;
        end
        else
        begin
          state       <=hb_dec_LdataB;
          memwra_en   <=(vncn_count==4'd4 | vncn_count==4'd6 | vncn_count==4'd8 | vncn_count==4'd10) ;
          memwrb_en   <=(ch_countb < 13'd656);
          if(layer_i==2'd3 & addr_count==4'd15 & vncn_count==4'd11 & section==2'd3)
            iter_count<=(iter_count==maxiter)?5'd8:iter_count +5'd1;
          if(addr_count==4'd15 & section==2'd3 & vncn_count==4'd11)
            layer_i   <=layer_i+2'd1;
          section     <=(vncn_count>=4'd4)? (~memwra_en)? section:section+2'd1:section+2'd1;
          addr_count  <=(section==2'd3 & vncn_count==4'd11)?addr_count+4'd1:addr_count;
          vncn_count  <=(vncn_count==4'd11)?4'd0:vncn_count+4'd1;
          hb_count    <=(hb_en)?(hb_count==4'd15)?4'd0:hb_count+4'd1:4'd0;
          dec_fin     <=0;
          hb_count_wr <=(section==2'd3 & vncn_count==4'd11)?hb_count_wr+4'd1:hb_count_wr;
          section_hb<=(hb_en)?((hb_count==4'd15)?
                       section_hb+2'd1:section_hb):2'd0 ;
          if(hb_vlid)
          begin
            if((hb_count==4'd0) & section_hb==2'd0)
              memid_hb<=(memid_hb==6'd15)? 6'd0 :
                     (~data_wrsa & ~data_wrsb)? 6'd0 : memid_hb+6'd1;
            if((memid_hb==6'd1 | memid_hb==6'd3 | memid_hb==6'd5 | memid_hb==6'd7 | memid_hb==6'd9) & (hb_count==4'd0) & section_hb==2'd0)
              memgroup_hb<=(memgroup_hb==3'd4)?
                         3'd0 : memgroup_hb+3'd1;
          end
        end
      end
      hb_act://state:4'b0111
      begin
        data_wrsa   <=0;
        data_wrsb   <=0;
        hb_vlid     <=(ch_counta >=13'd16 & ch_counta <13'd657);
        hb_en       <=1;
        load_data_en<=0;
        memwra_en   <=0;
        memwrb_en   <=0;
        ch_counta   <=(ch_counta==maxiter*768)?13'd0:ch_counta+13'd1;
        ch_countb   <=0;
        vncn_count  <=0;
        layer_i     <=0;
        section     <=0;
        addr_count  <=0;
        addr_ch_count<=0;
        iter_count  <=0;
        state       <=(~hb_vlid)?3'b010:hb_act;
        hb_count    <=(hb_en)?(hb_count==4'd15)?4'd0:hb_count+4'd1:4'd0;
        dec_fin     <=1;
        hb_count_wr <=0;
        memid_hb    <=0;
        memgroup_hb <=0;
        section_hb  <=0;
      end
      default:
      begin
        load_data_en<=0;
        memwra_en   <=0;
        memwrb_en   <=0;
        vncn_count  <=0;
        addr_count  <=0;
        addr_ch_count<=0;
        ch_counta   <=0;
        ch_countb   <=0;
        hb_count    <=0;
        layer_i     <=0;
        section     <=0;
        iter_count  <=0;
        hb_vlid     <=0;
        hb_en       <=0;
        data_wrsa   <=0;
        data_wrsb   <=0;
        state       <=(start_ldpc)?load_data:idle;
        dec_fin     <=1;
        hb_count_wr <=0;
        memid_hb    <=0;
        memgroup_hb <=0;
        section_hb  <=0;
      end
    endcase
  end
end
endmodule
module CMPtop(
           vtc_1,vtc_2,vtc_3,vtc_4,vtc_5,
           min,secmin,
           minaddr);

input  [1:0] vtc_1,vtc_2,vtc_3,vtc_4,vtc_5;
output [1:0] min,secmin;
output [4:0] minaddr;
wire   [1:0] min_tmp1,secmin_tmp1,min_tmp2,secmin_tmp2,min_tmp3,secmin_tmp3,min,secmin;
wire   [4:0] minaddr_tmp1,minaddr_tmp2,minaddr_tmp3,minaddr;

assign min_tmp1=(vtc_1>vtc_2)?vtc_2:vtc_1;
assign secmin_tmp1=(vtc_1>vtc_2)?vtc_1:vtc_2;
assign minaddr_tmp1=(vtc_1>vtc_2)?5'd2:5'd1;

assign min_tmp2=(min_tmp1 >vtc_3)?vtc_3:min_tmp1;
assign secmin_tmp2=(min_tmp1 >vtc_3)?min_tmp1:((secmin_tmp1>vtc_3) & (vtc_3!=min_tmp1))?vtc_3:secmin_tmp1;
assign minaddr_tmp2=(min_tmp1 >vtc_3)?5'd4:minaddr_tmp1;

assign min_tmp3=(min_tmp2 >vtc_4)?vtc_4:min_tmp2;
assign secmin_tmp3=(min_tmp2 >vtc_4)?min_tmp2:((secmin_tmp2>vtc_4) & (vtc_4!=min_tmp2))?vtc_4:secmin_tmp2;
assign minaddr_tmp3=(min_tmp2 >vtc_4)?5'd8:minaddr_tmp2;

assign min=(min_tmp3 >vtc_5)?vtc_5:min_tmp3;
assign secmin=(min_tmp3 >vtc_5)?min_tmp3:((secmin_tmp3>vtc_5) & (vtc_5!=min_tmp3))?vtc_5:secmin_tmp3;
assign minaddr=(min_tmp3 >vtc_5)?5'd16:minaddr_tmp3;
endmodule

module CNP(
           CLK,RESET_N,
           vncn_en,totsgn,keep_min,
           vtc_1,vtc_2,
           min_r,secmin_r,section,
           min_loc,
           ctm_1,ctm_2,
           min,
           sgn);

input        CLK,RESET_N;
input        vncn_en,totsgn,keep_min;
input  [2:0] vtc_1,vtc_2;
input  [1:0] min_r,secmin_r,section;
input        min_loc;
output [2:0] ctm_1,ctm_2;
output [1:0] min;
output sgn;

reg  [1:0] min;
reg  [2:0] minaddr; //rm1 for vncn rm2 for mem

reg [7:0] sgn_r;

wire [1:0]vtc1=(vtc_1[2])? (vtc_1[1] | vtc_1[0])?~vtc_1[1:0]+2'd1:2'b11:vtc_1[1:0];
wire [1:0]vtc2=(vtc_2[2])? (vtc_2[1] | vtc_2[0])?~vtc_2[1:0]+2'd1:2'b11:vtc_2[1:0];

wire [1:0] min1=(vtc1>vtc2)?vtc2:vtc1;
wire [2:0] minaddr1=(vtc1>vtc2)?3'd1:3'd0;
wire sgn=^sgn_r;
always @(negedge RESET_N or posedge CLK)
begin
  if (~RESET_N)
  begin
    min      <=2'd3;
    minaddr  <=0;
    sgn_r    <=0;
  end
  else if(vncn_en)
  begin
    min      <=2'd3;
    minaddr  <=0;
    sgn_r    <=0;
  end
  else if(~keep_min)
  begin
    if(min1<=min) min<=min1 ;
    if(min1<=min) minaddr<=minaddr1+{1'd0,section}+{1'd0,section};
    sgn_r<={vtc_1[2],vtc_2[2],sgn_r[7:2]};
  end
end

wire sgn1=(section==2'd0) ? sgn_r[1] :
          (section==2'd1) ? sgn_r[3] :
          (section==2'd2) ? sgn_r[5] : sgn_r[7];
  wire sgn2=(section==2'd0) ? sgn_r[0] :
          (section==2'd1) ? sgn_r[2] :
          (section==2'd2) ? sgn_r[4] : sgn_r[6];

wire [1:0] minsel1= ((section==2'd0 & minaddr==3'd0)|
                     (section==2'd1 & minaddr==3'd2)|
                     (section==2'd2 & minaddr==3'd4)|
                     (section==2'd3 & minaddr==3'd6)& min_loc)?
                      (secmin_r==2'd0)? 2'd0:secmin_r-2'd1 : (min_r==2'd0)? 2'd0:min_r-2'd1;
wire [1:0] minsel2= ((section==2'd0 & minaddr==3'd1)|
                     (section==2'd1 & minaddr==3'd3)|
                     (section==2'd2 & minaddr==3'd5)|
                     (section==2'd3 & minaddr==3'd7)& min_loc)?
                      (secmin_r==2'd0)? 2'd0:secmin_r-2'd1 : (min_r==2'd0)? 2'd0:min_r-2'd1;

wire [2:0] ctm_1=(totsgn^sgn1)?{totsgn^sgn1,~minsel1+2'd1}:{totsgn^sgn1,minsel1};
wire [2:0] ctm_2=(totsgn^sgn2)?{totsgn^sgn2,~minsel2+2'd1}:{totsgn^sgn2,minsel2};

endmodule

module memblock64x32(
            A,
            CEN,
            CLK,
            D,
            WEN,
            Q
                   );
input [5:0] A;
input CEN,CLK,WEN;
input [31:0] D;
output [31:0] Q;
reg [31:0] D_r [0:63];
reg [31:0] Q;
always @(posedge CLK)
if(WEN & CEN)
begin
  D_r[A]<=D;
  Q<=D_r[A];
end
else
begin
  Q<=D_r[A];
end
endmodule

module memblock256x48(
                      A,
                      CEN,
                      CLK,
                      D,
                      WEN,
                      Q
                      );
input [7:0] A;
input CEN,CLK,WEN;
input [47:0] D;
output [47:0] Q;
reg [47:0] D_r [0:255];
reg [47:0] Q;
always @(posedge CLK)
if(WEN & CEN)
begin
  D_r[A]<=D;
  Q<=D_r[A];
end
else
begin
  Q<=D_r[A];
end
endmodule

module memblock64x80(
                    A,
                    CEN,
                    CLK,
                    D,
                    WEN,
                    Q
                      );
input [5:0] A;
input CEN,CLK,WEN;
input [79:0] D;
output [79:0] Q;
reg [79:0] D_r [0:63];
reg [79:0] Q;
always @(posedge CLK)
if(WEN & CEN)
begin
  D_r[A]<=D;
  Q<=D_r[A];
end
else
begin
  Q<=D_r[A];
end
endmodule

                                 